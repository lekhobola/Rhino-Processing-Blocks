--********************************************************************************
--* Company:        University of Cape Town									   
--* Engineer:       Lekhobola Joachim Tsoeunyane, lekhobola@gmail.com		       
--********************************************************************************
--* Create Date:    06-Jul-2014 01:03:44  				 										   
--* Design Name:    Pipelined R2^2 DIF-SDF FFT								       
--* Module Name:    fft4096_tf_rom_s0.vhd										   
--* Project Name:   RHINO SDR Processing Blocks								   
--* Target Devices: Xilinx - SPARTAN-6											   
--********************************************************************************
--* Dependencies: none															   
--********************************************************************************
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--********************************************************************************
--* This module implements the stage-0 of twiddle factor ROM for a 4096-point      
--* pipelined R2^2 DIF-SDF FFT. Each value is a complex number{imaginary,complex} 
--* ******************************************************************************
--* params:																	   
--*        addr_w - rom address bit width									       
--*        data_w - output data bit width										   
--* ports:																		   
--* 			[in]  addr	- Twidde factor ROM address to read					   
--* 			[out] doutr - Twiddle factor read from rom addr - real value	   
--* 			[out] douti - Twidder factor read from rom addr - imaginary value  
--********************************************************************************
--* Notes: Do not modify this file as it is auto-generated using matlab script    
--********************************************************************************
entity fft4096_tf_rom_s0 is
	generic(
		addr_w : natural := 12;
		data_w : natural := 16
	);
    port (
        addr  : in  std_logic_vector (addr_w - 1 downto 0);
        doutr : out std_logic_vector (data_w - 1 downto 0);
        douti : out  std_logic_vector(data_w - 1 downto 0)
 	);
end fft4096_tf_rom_s0;

architecture Behavioral of fft4096_tf_rom_s0 is
	type complex is array(0 to 1) of std_logic_vector(data_w - 1 downto 0);
	type rom_type is array(0 to (2 ** addr_w) - 1) of complex;

	constant rom : rom_type := (
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","1111111111001110"),
								 ("0100000000000000","1111111110011011"),
								 ("0011111111111111","1111111101101001"),
								 ("0011111111111111","1111111100110111"),
								 ("0011111111111110","1111111100000101"),
								 ("0011111111111101","1111111011010010"),
								 ("0011111111111100","1111111010100000"),
								 ("0011111111111011","1111111001101110"),
								 ("0011111111111010","1111111000111100"),
								 ("0011111111111000","1111111000001001"),
								 ("0011111111110111","1111110111010111"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111110011","1111110101110011"),
								 ("0011111111110001","1111110101000000"),
								 ("0011111111101111","1111110100001110"),
								 ("0011111111101100","1111110011011100"),
								 ("0011111111101010","1111110010101010"),
								 ("0011111111100111","1111110001111000"),
								 ("0011111111100100","1111110001000101"),
								 ("0011111111100001","1111110000010011"),
								 ("0011111111011110","1111101111100001"),
								 ("0011111111011011","1111101110101111"),
								 ("0011111111010111","1111101101111101"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111111010000","1111101100011001"),
								 ("0011111111001100","1111101011100110"),
								 ("0011111111001000","1111101010110100"),
								 ("0011111111000100","1111101010000010"),
								 ("0011111110111111","1111101001010000"),
								 ("0011111110111011","1111101000011110"),
								 ("0011111110110110","1111100111101100"),
								 ("0011111110110001","1111100110111010"),
								 ("0011111110101100","1111100110001000"),
								 ("0011111110100111","1111100101010110"),
								 ("0011111110100010","1111100100100100"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111110010111","1111100011000000"),
								 ("0011111110010001","1111100010001110"),
								 ("0011111110001011","1111100001011100"),
								 ("0011111110000101","1111100000101010"),
								 ("0011111101111111","1111011111111001"),
								 ("0011111101111000","1111011111000111"),
								 ("0011111101110010","1111011110010101"),
								 ("0011111101101011","1111011101100011"),
								 ("0011111101100100","1111011100110001"),
								 ("0011111101011101","1111011011111111"),
								 ("0011111101010110","1111011011001110"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111101000111","1111011001101010"),
								 ("0011111101000000","1111011000111001"),
								 ("0011111100111000","1111011000000111"),
								 ("0011111100110000","1111010111010101"),
								 ("0011111100101000","1111010110100100"),
								 ("0011111100100000","1111010101110010"),
								 ("0011111100010111","1111010101000000"),
								 ("0011111100001111","1111010100001111"),
								 ("0011111100000110","1111010011011101"),
								 ("0011111011111101","1111010010101100"),
								 ("0011111011110100","1111010001111011"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111011100010","1111010000011000"),
								 ("0011111011011000","1111001111100110"),
								 ("0011111011001111","1111001110110101"),
								 ("0011111011000101","1111001110000100"),
								 ("0011111010111011","1111001101010010"),
								 ("0011111010110001","1111001100100001"),
								 ("0011111010100111","1111001011110000"),
								 ("0011111010011101","1111001010111111"),
								 ("0011111010010010","1111001010001110"),
								 ("0011111010001000","1111001001011100"),
								 ("0011111001111101","1111001000101011"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111001100111","1111000111001001"),
								 ("0011111001011100","1111000110011000"),
								 ("0011111001010000","1111000101100111"),
								 ("0011111001000101","1111000100110110"),
								 ("0011111000111001","1111000100000101"),
								 ("0011111000101101","1111000011010101"),
								 ("0011111000100001","1111000010100100"),
								 ("0011111000010101","1111000001110011"),
								 ("0011111000001001","1111000001000010"),
								 ("0011110111111100","1111000000010010"),
								 ("0011110111110000","1110111111100001"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110111010110","1110111110000000"),
								 ("0011110111001001","1110111101001111"),
								 ("0011110110111100","1110111100011111"),
								 ("0011110110101111","1110111011101110"),
								 ("0011110110100001","1110111010111110"),
								 ("0011110110010011","1110111010001101"),
								 ("0011110110000110","1110111001011101"),
								 ("0011110101111000","1110111000101101"),
								 ("0011110101101010","1110110111111100"),
								 ("0011110101011011","1110110111001100"),
								 ("0011110101001101","1110110110011100"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110100110000","1110110100111100"),
								 ("0011110100100001","1110110100001100"),
								 ("0011110100010010","1110110011011100"),
								 ("0011110100000011","1110110010101100"),
								 ("0011110011110100","1110110001111100"),
								 ("0011110011100100","1110110001001100"),
								 ("0011110011010101","1110110000011100"),
								 ("0011110011000101","1110101111101101"),
								 ("0011110010110101","1110101110111101"),
								 ("0011110010100101","1110101110001101"),
								 ("0011110010010101","1110101101011110"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110001110100","1110101011111111"),
								 ("0011110001100100","1110101011001111"),
								 ("0011110001010011","1110101010100000"),
								 ("0011110001000010","1110101001110000"),
								 ("0011110000110001","1110101001000001"),
								 ("0011110000100000","1110101000010010"),
								 ("0011110000001111","1110100111100011"),
								 ("0011101111111101","1110100110110100"),
								 ("0011101111101100","1110100110000100"),
								 ("0011101111011010","1110100101010101"),
								 ("0011101111001000","1110100100100110"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101110100100","1110100011001001"),
								 ("0011101110010010","1110100010011010"),
								 ("0011101101111111","1110100001101011"),
								 ("0011101101101101","1110100000111100"),
								 ("0011101101011010","1110100000001110"),
								 ("0011101101000111","1110011111011111"),
								 ("0011101100110100","1110011110110001"),
								 ("0011101100100001","1110011110000010"),
								 ("0011101100001110","1110011101010100"),
								 ("0011101011111010","1110011100100101"),
								 ("0011101011100110","1110011011110111"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101010111111","1110011010011011"),
								 ("0011101010101011","1110011001101101"),
								 ("0011101010010111","1110011000111111"),
								 ("0011101010000010","1110011000010001"),
								 ("0011101001101110","1110010111100011"),
								 ("0011101001011001","1110010110110101"),
								 ("0011101001000101","1110010110000111"),
								 ("0011101000110000","1110010101011001"),
								 ("0011101000011011","1110010100101100"),
								 ("0011101000000110","1110010011111110"),
								 ("0011100111110000","1110010011010000"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100111000101","1110010001110110"),
								 ("0011100110110000","1110010001001000"),
								 ("0011100110011010","1110010000011011"),
								 ("0011100110000100","1110001111101110"),
								 ("0011100101101110","1110001111000001"),
								 ("0011100101011000","1110001110010100"),
								 ("0011100101000001","1110001101100111"),
								 ("0011100100101011","1110001100111010"),
								 ("0011100100010100","1110001100001101"),
								 ("0011100011111101","1110001011100000"),
								 ("0011100011100110","1110001010110011"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100010111000","1110001001011010"),
								 ("0011100010100001","1110001000101101"),
								 ("0011100010001001","1110001000000001"),
								 ("0011100001110001","1110000111010101"),
								 ("0011100001011010","1110000110101000"),
								 ("0011100001000010","1110000101111100"),
								 ("0011100000101010","1110000101010000"),
								 ("0011100000010010","1110000100100100"),
								 ("0011011111111001","1110000011111000"),
								 ("0011011111100001","1110000011001100"),
								 ("0011011111001000","1110000010100000"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011110010111","1110000001001001"),
								 ("0011011101111110","1110000000011101"),
								 ("0011011101100101","1101111111110001"),
								 ("0011011101001011","1101111111000110"),
								 ("0011011100110010","1101111110011011"),
								 ("0011011100011000","1101111101101111"),
								 ("0011011011111111","1101111101000100"),
								 ("0011011011100101","1101111100011001"),
								 ("0011011011001011","1101111011101110"),
								 ("0011011010110001","1101111011000011"),
								 ("0011011010010111","1101111010011000"),
								 ("0011011001111101","1101111001101101"),
								 ("0011011001100010","1101111001000010"),
								 ("0011011001001000","1101111000011000"),
								 ("0011011000101101","1101110111101101"),
								 ("0011011000010010","1101110111000011"),
								 ("0011010111110111","1101110110011000"),
								 ("0011010111011100","1101110101101110"),
								 ("0011010111000001","1101110101000100"),
								 ("0011010110100101","1101110100011001"),
								 ("0011010110001010","1101110011101111"),
								 ("0011010101101110","1101110011000101"),
								 ("0011010101010011","1101110010011011"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010100011011","1101110001001000"),
								 ("0011010011111111","1101110000011110"),
								 ("0011010011100010","1101101111110101"),
								 ("0011010011000110","1101101111001011"),
								 ("0011010010101010","1101101110100010"),
								 ("0011010010001101","1101101101111000"),
								 ("0011010001110000","1101101101001111"),
								 ("0011010001010011","1101101100100110"),
								 ("0011010000110110","1101101011111101"),
								 ("0011010000011001","1101101011010100"),
								 ("0011001111111100","1101101010101011"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001111000001","1101101001011010"),
								 ("0011001110100011","1101101000110001"),
								 ("0011001110000110","1101101000001000"),
								 ("0011001101101000","1101100111100000"),
								 ("0011001101001010","1101100110111000"),
								 ("0011001100101100","1101100110001111"),
								 ("0011001100001101","1101100101100111"),
								 ("0011001011101111","1101100100111111"),
								 ("0011001011010000","1101100100010111"),
								 ("0011001010110010","1101100011101111"),
								 ("0011001010010011","1101100011001000"),
								 ("0011001001110100","1101100010100000"),
								 ("0011001001010101","1101100001111000"),
								 ("0011001000110110","1101100001010001"),
								 ("0011001000010111","1101100000101010"),
								 ("0011000111111000","1101100000000010"),
								 ("0011000111011000","1101011111011011"),
								 ("0011000110111001","1101011110110100"),
								 ("0011000110011001","1101011110001101"),
								 ("0011000101111001","1101011101100110"),
								 ("0011000101011001","1101011100111111"),
								 ("0011000100111001","1101011100011001"),
								 ("0011000100011001","1101011011110010"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000011011000","1101011010100101"),
								 ("0011000010111000","1101011001111111"),
								 ("0011000010010111","1101011001011001"),
								 ("0011000001110110","1101011000110010"),
								 ("0011000001010101","1101011000001100"),
								 ("0011000000110100","1101010111100110"),
								 ("0011000000010011","1101010111000001"),
								 ("0010111111110010","1101010110011011"),
								 ("0010111111010000","1101010101110101"),
								 ("0010111110101111","1101010101010000"),
								 ("0010111110001101","1101010100101010"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111101001010","1101010011100000"),
								 ("0010111100101000","1101010010111011"),
								 ("0010111100000110","1101010010010110"),
								 ("0010111011100100","1101010001110001"),
								 ("0010111011000010","1101010001001100"),
								 ("0010111010011111","1101010000101000"),
								 ("0010111001111101","1101010000000011"),
								 ("0010111001011010","1101001111011111"),
								 ("0010111000110111","1101001110111010"),
								 ("0010111000010101","1101001110010110"),
								 ("0010110111110010","1101001101110010"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110110101011","1101001100101010"),
								 ("0010110110001000","1101001100000110"),
								 ("0010110101100101","1101001011100010"),
								 ("0010110101000001","1101001010111111"),
								 ("0010110100011110","1101001010011011"),
								 ("0010110011111010","1101001001111000"),
								 ("0010110011010110","1101001001010101"),
								 ("0010110010110010","1101001000110001"),
								 ("0010110010001110","1101001000001110"),
								 ("0010110001101010","1101000111101011"),
								 ("0010110001000110","1101000111001001"),
								 ("0010110000100001","1101000110100110"),
								 ("0010101111111101","1101000110000011"),
								 ("0010101111011000","1101000101100001"),
								 ("0010101110110100","1101000100111110"),
								 ("0010101110001111","1101000100011100"),
								 ("0010101101101010","1101000011111010"),
								 ("0010101101000101","1101000011011000"),
								 ("0010101100100000","1101000010110110"),
								 ("0010101011111011","1101000010010100"),
								 ("0010101011010110","1101000001110011"),
								 ("0010101010110000","1101000001010001"),
								 ("0010101010001011","1101000000110000"),
								 ("0010101001100101","1101000000001110"),
								 ("0010101000111111","1100111111101101"),
								 ("0010101000011010","1100111111001100"),
								 ("0010100111110100","1100111110101011"),
								 ("0010100111001110","1100111110001010"),
								 ("0010100110100111","1100111101101001"),
								 ("0010100110000001","1100111101001000"),
								 ("0010100101011011","1100111100101000"),
								 ("0010100100110101","1100111100000111"),
								 ("0010100100001110","1100111011100111"),
								 ("0010100011100111","1100111011000111"),
								 ("0010100011000001","1100111010100111"),
								 ("0010100010011010","1100111010000111"),
								 ("0010100001110011","1100111001100111"),
								 ("0010100001001100","1100111001000111"),
								 ("0010100000100101","1100111000101000"),
								 ("0010011111111110","1100111000001000"),
								 ("0010011111010110","1100110111101001"),
								 ("0010011110101111","1100110111001010"),
								 ("0010011110001000","1100110110101011"),
								 ("0010011101100000","1100110110001100"),
								 ("0010011100111000","1100110101101101"),
								 ("0010011100010001","1100110101001110"),
								 ("0010011011101001","1100110100110000"),
								 ("0010011011000001","1100110100010001"),
								 ("0010011010011001","1100110011110011"),
								 ("0010011001110001","1100110011010100"),
								 ("0010011001001000","1100110010110110"),
								 ("0010011000100000","1100110010011000"),
								 ("0010010111111000","1100110001111010"),
								 ("0010010111001111","1100110001011101"),
								 ("0010010110100110","1100110000111111"),
								 ("0010010101111110","1100110000100001"),
								 ("0010010101010101","1100110000000100"),
								 ("0010010100101100","1100101111100111"),
								 ("0010010100000011","1100101111001010"),
								 ("0010010011011010","1100101110101101"),
								 ("0010010010110001","1100101110010000"),
								 ("0010010010001000","1100101101110011"),
								 ("0010010001011110","1100101101010110"),
								 ("0010010000110101","1100101100111010"),
								 ("0010010000001011","1100101100011110"),
								 ("0010001111100010","1100101100000001"),
								 ("0010001110111000","1100101011100101"),
								 ("0010001110001110","1100101011001001"),
								 ("0010001101100101","1100101010101101"),
								 ("0010001100111011","1100101010010010"),
								 ("0010001100010001","1100101001110110"),
								 ("0010001011100111","1100101001011011"),
								 ("0010001010111100","1100101000111111"),
								 ("0010001010010010","1100101000100100"),
								 ("0010001001101000","1100101000001001"),
								 ("0010001000111101","1100100111101110"),
								 ("0010001000010011","1100100111010011"),
								 ("0010000111101000","1100100110111000"),
								 ("0010000110111110","1100100110011110"),
								 ("0010000110010011","1100100110000011"),
								 ("0010000101101000","1100100101101001"),
								 ("0010000100111101","1100100101001111"),
								 ("0010000100010010","1100100100110101"),
								 ("0010000011100111","1100100100011011"),
								 ("0010000010111100","1100100100000001"),
								 ("0010000010010001","1100100011101000"),
								 ("0010000001100101","1100100011001110"),
								 ("0010000000111010","1100100010110101"),
								 ("0010000000001111","1100100010011011"),
								 ("0001111111100011","1100100010000010"),
								 ("0001111110110111","1100100001101001"),
								 ("0001111110001100","1100100001010000"),
								 ("0001111101100000","1100100000111000"),
								 ("0001111100110100","1100100000011111"),
								 ("0001111100001000","1100100000000111"),
								 ("0001111011011100","1100011111101110"),
								 ("0001111010110000","1100011111010110"),
								 ("0001111010000100","1100011110111110"),
								 ("0001111001011000","1100011110100110"),
								 ("0001111000101011","1100011110001111"),
								 ("0001110111111111","1100011101110111"),
								 ("0001110111010011","1100011101011111"),
								 ("0001110110100110","1100011101001000"),
								 ("0001110101111001","1100011100110001"),
								 ("0001110101001101","1100011100011010"),
								 ("0001110100100000","1100011100000011"),
								 ("0001110011110011","1100011011101100"),
								 ("0001110011000110","1100011011010101"),
								 ("0001110010011001","1100011010111111"),
								 ("0001110001101100","1100011010101000"),
								 ("0001110000111111","1100011010010010"),
								 ("0001110000010010","1100011001111100"),
								 ("0001101111100101","1100011001100110"),
								 ("0001101110111000","1100011001010000"),
								 ("0001101110001010","1100011000111011"),
								 ("0001101101011101","1100011000100101"),
								 ("0001101100110000","1100011000010000"),
								 ("0001101100000010","1100010111111010"),
								 ("0001101011010100","1100010111100101"),
								 ("0001101010100111","1100010111010000"),
								 ("0001101001111001","1100010110111011"),
								 ("0001101001001011","1100010110100111"),
								 ("0001101000011101","1100010110010010"),
								 ("0001100111101111","1100010101111110"),
								 ("0001100111000001","1100010101101001"),
								 ("0001100110010011","1100010101010101"),
								 ("0001100101100101","1100010101000001"),
								 ("0001100100110111","1100010100101101"),
								 ("0001100100001001","1100010100011010"),
								 ("0001100011011011","1100010100000110"),
								 ("0001100010101100","1100010011110010"),
								 ("0001100001111110","1100010011011111"),
								 ("0001100001001111","1100010011001100"),
								 ("0001100000100001","1100010010111001"),
								 ("0001011111110010","1100010010100110"),
								 ("0001011111000100","1100010010010011"),
								 ("0001011110010101","1100010010000001"),
								 ("0001011101100110","1100010001101110"),
								 ("0001011100110111","1100010001011100"),
								 ("0001011100001001","1100010001001010"),
								 ("0001011011011010","1100010000111000"),
								 ("0001011010101011","1100010000100110"),
								 ("0001011001111100","1100010000010100"),
								 ("0001011001001100","1100010000000011"),
								 ("0001011000011101","1100001111110001"),
								 ("0001010111101110","1100001111100000"),
								 ("0001010110111111","1100001111001111"),
								 ("0001010110010000","1100001110111110"),
								 ("0001010101100000","1100001110101101"),
								 ("0001010100110001","1100001110011100"),
								 ("0001010100000001","1100001110001100"),
								 ("0001010011010010","1100001101111011"),
								 ("0001010010100010","1100001101101011"),
								 ("0001010001110011","1100001101011011"),
								 ("0001010001000011","1100001101001011"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001111100100","1100001100101011"),
								 ("0001001110110100","1100001100011100"),
								 ("0001001110000100","1100001100001100"),
								 ("0001001101010100","1100001011111101"),
								 ("0001001100100100","1100001011101110"),
								 ("0001001011110100","1100001011011111"),
								 ("0001001011000100","1100001011010000"),
								 ("0001001010010100","1100001011000001"),
								 ("0001001001100100","1100001010110011"),
								 ("0001001000110100","1100001010100101"),
								 ("0001001000000100","1100001010010110"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000110100011","1100001001111010"),
								 ("0001000101110011","1100001001101101"),
								 ("0001000101000010","1100001001011111"),
								 ("0001000100010010","1100001001010001"),
								 ("0001000011100001","1100001001000100"),
								 ("0001000010110001","1100001000110111"),
								 ("0001000010000000","1100001000101010"),
								 ("0001000001010000","1100001000011101"),
								 ("0001000000011111","1100001000010000"),
								 ("0000111111101110","1100001000000100"),
								 ("0000111110111110","1100000111110111"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111101011100","1100000111011111"),
								 ("0000111100101011","1100000111010011"),
								 ("0000111011111011","1100000111000111"),
								 ("0000111011001010","1100000110111011"),
								 ("0000111010011001","1100000110110000"),
								 ("0000111001101000","1100000110100100"),
								 ("0000111000110111","1100000110011001"),
								 ("0000111000000110","1100000110001110"),
								 ("0000110111010101","1100000110000011"),
								 ("0000110110100100","1100000101111000"),
								 ("0000110101110010","1100000101101110"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110100010000","1100000101011001"),
								 ("0000110011011111","1100000101001111"),
								 ("0000110010101110","1100000101000101"),
								 ("0000110001111100","1100000100111011"),
								 ("0000110001001011","1100000100110001"),
								 ("0000110000011010","1100000100101000"),
								 ("0000101111101000","1100000100011110"),
								 ("0000101110110111","1100000100010101"),
								 ("0000101110000101","1100000100001100"),
								 ("0000101101010100","1100000100000011"),
								 ("0000101100100011","1100000011111010"),
								 ("0000101011110001","1100000011110001"),
								 ("0000101011000000","1100000011101001"),
								 ("0000101010001110","1100000011100000"),
								 ("0000101001011100","1100000011011000"),
								 ("0000101000101011","1100000011010000"),
								 ("0000100111111001","1100000011001000"),
								 ("0000100111000111","1100000011000000"),
								 ("0000100110010110","1100000010111001"),
								 ("0000100101100100","1100000010110001"),
								 ("0000100100110010","1100000010101010"),
								 ("0000100100000001","1100000010100011"),
								 ("0000100011001111","1100000010011100"),
								 ("0000100010011101","1100000010010101"),
								 ("0000100001101011","1100000010001110"),
								 ("0000100000111001","1100000010001000"),
								 ("0000100000000111","1100000010000001"),
								 ("0000011111010110","1100000001111011"),
								 ("0000011110100100","1100000001110101"),
								 ("0000011101110010","1100000001101111"),
								 ("0000011101000000","1100000001101001"),
								 ("0000011100001110","1100000001100100"),
								 ("0000011011011100","1100000001011110"),
								 ("0000011010101010","1100000001011001"),
								 ("0000011001111000","1100000001010100"),
								 ("0000011001000110","1100000001001111"),
								 ("0000011000010100","1100000001001010"),
								 ("0000010111100010","1100000001000101"),
								 ("0000010110110000","1100000001000001"),
								 ("0000010101111110","1100000000111100"),
								 ("0000010101001100","1100000000111000"),
								 ("0000010100011010","1100000000110100"),
								 ("0000010011100111","1100000000110000"),
								 ("0000010010110101","1100000000101100"),
								 ("0000010010000011","1100000000101001"),
								 ("0000010001010001","1100000000100101"),
								 ("0000010000011111","1100000000100010"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001110111011","1100000000011100"),
								 ("0000001110001000","1100000000011001"),
								 ("0000001101010110","1100000000010110"),
								 ("0000001100100100","1100000000010100"),
								 ("0000001011110010","1100000000010001"),
								 ("0000001011000000","1100000000001111"),
								 ("0000001010001101","1100000000001101"),
								 ("0000001001011011","1100000000001011"),
								 ("0000001000101001","1100000000001001"),
								 ("0000000111110111","1100000000001000"),
								 ("0000000111000100","1100000000000110"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000101100000","1100000000000100"),
								 ("0000000100101110","1100000000000011"),
								 ("0000000011111011","1100000000000010"),
								 ("0000000011001001","1100000000000001"),
								 ("0000000010010111","1100000000000001"),
								 ("0000000001100101","1100000000000000"),
								 ("0000000000110010","1100000000000000"),
								 ("0000000000000000","1100000000000000"),
								 ("1111111111001110","1100000000000000"),
								 ("1111111110011011","1100000000000000"),
								 ("1111111101101001","1100000000000001"),
								 ("1111111100110111","1100000000000001"),
								 ("1111111100000101","1100000000000010"),
								 ("1111111011010010","1100000000000011"),
								 ("1111111010100000","1100000000000100"),
								 ("1111111001101110","1100000000000101"),
								 ("1111111000111100","1100000000000110"),
								 ("1111111000001001","1100000000001000"),
								 ("1111110111010111","1100000000001001"),
								 ("1111110110100101","1100000000001011"),
								 ("1111110101110011","1100000000001101"),
								 ("1111110101000000","1100000000001111"),
								 ("1111110100001110","1100000000010001"),
								 ("1111110011011100","1100000000010100"),
								 ("1111110010101010","1100000000010110"),
								 ("1111110001111000","1100000000011001"),
								 ("1111110001000101","1100000000011100"),
								 ("1111110000010011","1100000000011111"),
								 ("1111101111100001","1100000000100010"),
								 ("1111101110101111","1100000000100101"),
								 ("1111101101111101","1100000000101001"),
								 ("1111101101001011","1100000000101100"),
								 ("1111101100011001","1100000000110000"),
								 ("1111101011100110","1100000000110100"),
								 ("1111101010110100","1100000000111000"),
								 ("1111101010000010","1100000000111100"),
								 ("1111101001010000","1100000001000001"),
								 ("1111101000011110","1100000001000101"),
								 ("1111100111101100","1100000001001010"),
								 ("1111100110111010","1100000001001111"),
								 ("1111100110001000","1100000001010100"),
								 ("1111100101010110","1100000001011001"),
								 ("1111100100100100","1100000001011110"),
								 ("1111100011110010","1100000001100100"),
								 ("1111100011000000","1100000001101001"),
								 ("1111100010001110","1100000001101111"),
								 ("1111100001011100","1100000001110101"),
								 ("1111100000101010","1100000001111011"),
								 ("1111011111111001","1100000010000001"),
								 ("1111011111000111","1100000010001000"),
								 ("1111011110010101","1100000010001110"),
								 ("1111011101100011","1100000010010101"),
								 ("1111011100110001","1100000010011100"),
								 ("1111011011111111","1100000010100011"),
								 ("1111011011001110","1100000010101010"),
								 ("1111011010011100","1100000010110001"),
								 ("1111011001101010","1100000010111001"),
								 ("1111011000111001","1100000011000000"),
								 ("1111011000000111","1100000011001000"),
								 ("1111010111010101","1100000011010000"),
								 ("1111010110100100","1100000011011000"),
								 ("1111010101110010","1100000011100000"),
								 ("1111010101000000","1100000011101001"),
								 ("1111010100001111","1100000011110001"),
								 ("1111010011011101","1100000011111010"),
								 ("1111010010101100","1100000100000011"),
								 ("1111010001111011","1100000100001100"),
								 ("1111010001001001","1100000100010101"),
								 ("1111010000011000","1100000100011110"),
								 ("1111001111100110","1100000100101000"),
								 ("1111001110110101","1100000100110001"),
								 ("1111001110000100","1100000100111011"),
								 ("1111001101010010","1100000101000101"),
								 ("1111001100100001","1100000101001111"),
								 ("1111001011110000","1100000101011001"),
								 ("1111001010111111","1100000101100011"),
								 ("1111001010001110","1100000101101110"),
								 ("1111001001011100","1100000101111000"),
								 ("1111001000101011","1100000110000011"),
								 ("1111000111111010","1100000110001110"),
								 ("1111000111001001","1100000110011001"),
								 ("1111000110011000","1100000110100100"),
								 ("1111000101100111","1100000110110000"),
								 ("1111000100110110","1100000110111011"),
								 ("1111000100000101","1100000111000111"),
								 ("1111000011010101","1100000111010011"),
								 ("1111000010100100","1100000111011111"),
								 ("1111000001110011","1100000111101011"),
								 ("1111000001000010","1100000111110111"),
								 ("1111000000010010","1100001000000100"),
								 ("1110111111100001","1100001000010000"),
								 ("1110111110110000","1100001000011101"),
								 ("1110111110000000","1100001000101010"),
								 ("1110111101001111","1100001000110111"),
								 ("1110111100011111","1100001001000100"),
								 ("1110111011101110","1100001001010001"),
								 ("1110111010111110","1100001001011111"),
								 ("1110111010001101","1100001001101101"),
								 ("1110111001011101","1100001001111010"),
								 ("1110111000101101","1100001010001000"),
								 ("1110110111111100","1100001010010110"),
								 ("1110110111001100","1100001010100101"),
								 ("1110110110011100","1100001010110011"),
								 ("1110110101101100","1100001011000001"),
								 ("1110110100111100","1100001011010000"),
								 ("1110110100001100","1100001011011111"),
								 ("1110110011011100","1100001011101110"),
								 ("1110110010101100","1100001011111101"),
								 ("1110110001111100","1100001100001100"),
								 ("1110110001001100","1100001100011100"),
								 ("1110110000011100","1100001100101011"),
								 ("1110101111101101","1100001100111011"),
								 ("1110101110111101","1100001101001011"),
								 ("1110101110001101","1100001101011011"),
								 ("1110101101011110","1100001101101011"),
								 ("1110101100101110","1100001101111011"),
								 ("1110101011111111","1100001110001100"),
								 ("1110101011001111","1100001110011100"),
								 ("1110101010100000","1100001110101101"),
								 ("1110101001110000","1100001110111110"),
								 ("1110101001000001","1100001111001111"),
								 ("1110101000010010","1100001111100000"),
								 ("1110100111100011","1100001111110001"),
								 ("1110100110110100","1100010000000011"),
								 ("1110100110000100","1100010000010100"),
								 ("1110100101010101","1100010000100110"),
								 ("1110100100100110","1100010000111000"),
								 ("1110100011110111","1100010001001010"),
								 ("1110100011001001","1100010001011100"),
								 ("1110100010011010","1100010001101110"),
								 ("1110100001101011","1100010010000001"),
								 ("1110100000111100","1100010010010011"),
								 ("1110100000001110","1100010010100110"),
								 ("1110011111011111","1100010010111001"),
								 ("1110011110110001","1100010011001100"),
								 ("1110011110000010","1100010011011111"),
								 ("1110011101010100","1100010011110010"),
								 ("1110011100100101","1100010100000110"),
								 ("1110011011110111","1100010100011010"),
								 ("1110011011001001","1100010100101101"),
								 ("1110011010011011","1100010101000001"),
								 ("1110011001101101","1100010101010101"),
								 ("1110011000111111","1100010101101001"),
								 ("1110011000010001","1100010101111110"),
								 ("1110010111100011","1100010110010010"),
								 ("1110010110110101","1100010110100111"),
								 ("1110010110000111","1100010110111011"),
								 ("1110010101011001","1100010111010000"),
								 ("1110010100101100","1100010111100101"),
								 ("1110010011111110","1100010111111010"),
								 ("1110010011010000","1100011000010000"),
								 ("1110010010100011","1100011000100101"),
								 ("1110010001110110","1100011000111011"),
								 ("1110010001001000","1100011001010000"),
								 ("1110010000011011","1100011001100110"),
								 ("1110001111101110","1100011001111100"),
								 ("1110001111000001","1100011010010010"),
								 ("1110001110010100","1100011010101000"),
								 ("1110001101100111","1100011010111111"),
								 ("1110001100111010","1100011011010101"),
								 ("1110001100001101","1100011011101100"),
								 ("1110001011100000","1100011100000011"),
								 ("1110001010110011","1100011100011010"),
								 ("1110001010000111","1100011100110001"),
								 ("1110001001011010","1100011101001000"),
								 ("1110001000101101","1100011101011111"),
								 ("1110001000000001","1100011101110111"),
								 ("1110000111010101","1100011110001111"),
								 ("1110000110101000","1100011110100110"),
								 ("1110000101111100","1100011110111110"),
								 ("1110000101010000","1100011111010110"),
								 ("1110000100100100","1100011111101110"),
								 ("1110000011111000","1100100000000111"),
								 ("1110000011001100","1100100000011111"),
								 ("1110000010100000","1100100000111000"),
								 ("1110000001110100","1100100001010000"),
								 ("1110000001001001","1100100001101001"),
								 ("1110000000011101","1100100010000010"),
								 ("1101111111110001","1100100010011011"),
								 ("1101111111000110","1100100010110101"),
								 ("1101111110011011","1100100011001110"),
								 ("1101111101101111","1100100011101000"),
								 ("1101111101000100","1100100100000001"),
								 ("1101111100011001","1100100100011011"),
								 ("1101111011101110","1100100100110101"),
								 ("1101111011000011","1100100101001111"),
								 ("1101111010011000","1100100101101001"),
								 ("1101111001101101","1100100110000011"),
								 ("1101111001000010","1100100110011110"),
								 ("1101111000011000","1100100110111000"),
								 ("1101110111101101","1100100111010011"),
								 ("1101110111000011","1100100111101110"),
								 ("1101110110011000","1100101000001001"),
								 ("1101110101101110","1100101000100100"),
								 ("1101110101000100","1100101000111111"),
								 ("1101110100011001","1100101001011011"),
								 ("1101110011101111","1100101001110110"),
								 ("1101110011000101","1100101010010010"),
								 ("1101110010011011","1100101010101101"),
								 ("1101110001110010","1100101011001001"),
								 ("1101110001001000","1100101011100101"),
								 ("1101110000011110","1100101100000001"),
								 ("1101101111110101","1100101100011110"),
								 ("1101101111001011","1100101100111010"),
								 ("1101101110100010","1100101101010110"),
								 ("1101101101111000","1100101101110011"),
								 ("1101101101001111","1100101110010000"),
								 ("1101101100100110","1100101110101101"),
								 ("1101101011111101","1100101111001010"),
								 ("1101101011010100","1100101111100111"),
								 ("1101101010101011","1100110000000100"),
								 ("1101101010000010","1100110000100001"),
								 ("1101101001011010","1100110000111111"),
								 ("1101101000110001","1100110001011101"),
								 ("1101101000001000","1100110001111010"),
								 ("1101100111100000","1100110010011000"),
								 ("1101100110111000","1100110010110110"),
								 ("1101100110001111","1100110011010100"),
								 ("1101100101100111","1100110011110011"),
								 ("1101100100111111","1100110100010001"),
								 ("1101100100010111","1100110100110000"),
								 ("1101100011101111","1100110101001110"),
								 ("1101100011001000","1100110101101101"),
								 ("1101100010100000","1100110110001100"),
								 ("1101100001111000","1100110110101011"),
								 ("1101100001010001","1100110111001010"),
								 ("1101100000101010","1100110111101001"),
								 ("1101100000000010","1100111000001000"),
								 ("1101011111011011","1100111000101000"),
								 ("1101011110110100","1100111001000111"),
								 ("1101011110001101","1100111001100111"),
								 ("1101011101100110","1100111010000111"),
								 ("1101011100111111","1100111010100111"),
								 ("1101011100011001","1100111011000111"),
								 ("1101011011110010","1100111011100111"),
								 ("1101011011001011","1100111100000111"),
								 ("1101011010100101","1100111100101000"),
								 ("1101011001111111","1100111101001000"),
								 ("1101011001011001","1100111101101001"),
								 ("1101011000110010","1100111110001010"),
								 ("1101011000001100","1100111110101011"),
								 ("1101010111100110","1100111111001100"),
								 ("1101010111000001","1100111111101101"),
								 ("1101010110011011","1101000000001110"),
								 ("1101010101110101","1101000000110000"),
								 ("1101010101010000","1101000001010001"),
								 ("1101010100101010","1101000001110011"),
								 ("1101010100000101","1101000010010100"),
								 ("1101010011100000","1101000010110110"),
								 ("1101010010111011","1101000011011000"),
								 ("1101010010010110","1101000011111010"),
								 ("1101010001110001","1101000100011100"),
								 ("1101010001001100","1101000100111110"),
								 ("1101010000101000","1101000101100001"),
								 ("1101010000000011","1101000110000011"),
								 ("1101001111011111","1101000110100110"),
								 ("1101001110111010","1101000111001001"),
								 ("1101001110010110","1101000111101011"),
								 ("1101001101110010","1101001000001110"),
								 ("1101001101001110","1101001000110001"),
								 ("1101001100101010","1101001001010101"),
								 ("1101001100000110","1101001001111000"),
								 ("1101001011100010","1101001010011011"),
								 ("1101001010111111","1101001010111111"),
								 ("1101001010011011","1101001011100010"),
								 ("1101001001111000","1101001100000110"),
								 ("1101001001010101","1101001100101010"),
								 ("1101001000110001","1101001101001110"),
								 ("1101001000001110","1101001101110010"),
								 ("1101000111101011","1101001110010110"),
								 ("1101000111001001","1101001110111010"),
								 ("1101000110100110","1101001111011111"),
								 ("1101000110000011","1101010000000011"),
								 ("1101000101100001","1101010000101000"),
								 ("1101000100111110","1101010001001100"),
								 ("1101000100011100","1101010001110001"),
								 ("1101000011111010","1101010010010110"),
								 ("1101000011011000","1101010010111011"),
								 ("1101000010110110","1101010011100000"),
								 ("1101000010010100","1101010100000101"),
								 ("1101000001110011","1101010100101010"),
								 ("1101000001010001","1101010101010000"),
								 ("1101000000110000","1101010101110101"),
								 ("1101000000001110","1101010110011011"),
								 ("1100111111101101","1101010111000001"),
								 ("1100111111001100","1101010111100110"),
								 ("1100111110101011","1101011000001100"),
								 ("1100111110001010","1101011000110010"),
								 ("1100111101101001","1101011001011001"),
								 ("1100111101001000","1101011001111111"),
								 ("1100111100101000","1101011010100101"),
								 ("1100111100000111","1101011011001011"),
								 ("1100111011100111","1101011011110010"),
								 ("1100111011000111","1101011100011001"),
								 ("1100111010100111","1101011100111111"),
								 ("1100111010000111","1101011101100110"),
								 ("1100111001100111","1101011110001101"),
								 ("1100111001000111","1101011110110100"),
								 ("1100111000101000","1101011111011011"),
								 ("1100111000001000","1101100000000010"),
								 ("1100110111101001","1101100000101010"),
								 ("1100110111001010","1101100001010001"),
								 ("1100110110101011","1101100001111000"),
								 ("1100110110001100","1101100010100000"),
								 ("1100110101101101","1101100011001000"),
								 ("1100110101001110","1101100011101111"),
								 ("1100110100110000","1101100100010111"),
								 ("1100110100010001","1101100100111111"),
								 ("1100110011110011","1101100101100111"),
								 ("1100110011010100","1101100110001111"),
								 ("1100110010110110","1101100110111000"),
								 ("1100110010011000","1101100111100000"),
								 ("1100110001111010","1101101000001000"),
								 ("1100110001011101","1101101000110001"),
								 ("1100110000111111","1101101001011010"),
								 ("1100110000100001","1101101010000010"),
								 ("1100110000000100","1101101010101011"),
								 ("1100101111100111","1101101011010100"),
								 ("1100101111001010","1101101011111101"),
								 ("1100101110101101","1101101100100110"),
								 ("1100101110010000","1101101101001111"),
								 ("1100101101110011","1101101101111000"),
								 ("1100101101010110","1101101110100010"),
								 ("1100101100111010","1101101111001011"),
								 ("1100101100011110","1101101111110101"),
								 ("1100101100000001","1101110000011110"),
								 ("1100101011100101","1101110001001000"),
								 ("1100101011001001","1101110001110010"),
								 ("1100101010101101","1101110010011011"),
								 ("1100101010010010","1101110011000101"),
								 ("1100101001110110","1101110011101111"),
								 ("1100101001011011","1101110100011001"),
								 ("1100101000111111","1101110101000100"),
								 ("1100101000100100","1101110101101110"),
								 ("1100101000001001","1101110110011000"),
								 ("1100100111101110","1101110111000011"),
								 ("1100100111010011","1101110111101101"),
								 ("1100100110111000","1101111000011000"),
								 ("1100100110011110","1101111001000010"),
								 ("1100100110000011","1101111001101101"),
								 ("1100100101101001","1101111010011000"),
								 ("1100100101001111","1101111011000011"),
								 ("1100100100110101","1101111011101110"),
								 ("1100100100011011","1101111100011001"),
								 ("1100100100000001","1101111101000100"),
								 ("1100100011101000","1101111101101111"),
								 ("1100100011001110","1101111110011011"),
								 ("1100100010110101","1101111111000110"),
								 ("1100100010011011","1101111111110001"),
								 ("1100100010000010","1110000000011101"),
								 ("1100100001101001","1110000001001001"),
								 ("1100100001010000","1110000001110100"),
								 ("1100100000111000","1110000010100000"),
								 ("1100100000011111","1110000011001100"),
								 ("1100100000000111","1110000011111000"),
								 ("1100011111101110","1110000100100100"),
								 ("1100011111010110","1110000101010000"),
								 ("1100011110111110","1110000101111100"),
								 ("1100011110100110","1110000110101000"),
								 ("1100011110001111","1110000111010101"),
								 ("1100011101110111","1110001000000001"),
								 ("1100011101011111","1110001000101101"),
								 ("1100011101001000","1110001001011010"),
								 ("1100011100110001","1110001010000111"),
								 ("1100011100011010","1110001010110011"),
								 ("1100011100000011","1110001011100000"),
								 ("1100011011101100","1110001100001101"),
								 ("1100011011010101","1110001100111010"),
								 ("1100011010111111","1110001101100111"),
								 ("1100011010101000","1110001110010100"),
								 ("1100011010010010","1110001111000001"),
								 ("1100011001111100","1110001111101110"),
								 ("1100011001100110","1110010000011011"),
								 ("1100011001010000","1110010001001000"),
								 ("1100011000111011","1110010001110110"),
								 ("1100011000100101","1110010010100011"),
								 ("1100011000010000","1110010011010000"),
								 ("1100010111111010","1110010011111110"),
								 ("1100010111100101","1110010100101100"),
								 ("1100010111010000","1110010101011001"),
								 ("1100010110111011","1110010110000111"),
								 ("1100010110100111","1110010110110101"),
								 ("1100010110010010","1110010111100011"),
								 ("1100010101111110","1110011000010001"),
								 ("1100010101101001","1110011000111111"),
								 ("1100010101010101","1110011001101101"),
								 ("1100010101000001","1110011010011011"),
								 ("1100010100101101","1110011011001001"),
								 ("1100010100011010","1110011011110111"),
								 ("1100010100000110","1110011100100101"),
								 ("1100010011110010","1110011101010100"),
								 ("1100010011011111","1110011110000010"),
								 ("1100010011001100","1110011110110001"),
								 ("1100010010111001","1110011111011111"),
								 ("1100010010100110","1110100000001110"),
								 ("1100010010010011","1110100000111100"),
								 ("1100010010000001","1110100001101011"),
								 ("1100010001101110","1110100010011010"),
								 ("1100010001011100","1110100011001001"),
								 ("1100010001001010","1110100011110111"),
								 ("1100010000111000","1110100100100110"),
								 ("1100010000100110","1110100101010101"),
								 ("1100010000010100","1110100110000100"),
								 ("1100010000000011","1110100110110100"),
								 ("1100001111110001","1110100111100011"),
								 ("1100001111100000","1110101000010010"),
								 ("1100001111001111","1110101001000001"),
								 ("1100001110111110","1110101001110000"),
								 ("1100001110101101","1110101010100000"),
								 ("1100001110011100","1110101011001111"),
								 ("1100001110001100","1110101011111111"),
								 ("1100001101111011","1110101100101110"),
								 ("1100001101101011","1110101101011110"),
								 ("1100001101011011","1110101110001101"),
								 ("1100001101001011","1110101110111101"),
								 ("1100001100111011","1110101111101101"),
								 ("1100001100101011","1110110000011100"),
								 ("1100001100011100","1110110001001100"),
								 ("1100001100001100","1110110001111100"),
								 ("1100001011111101","1110110010101100"),
								 ("1100001011101110","1110110011011100"),
								 ("1100001011011111","1110110100001100"),
								 ("1100001011010000","1110110100111100"),
								 ("1100001011000001","1110110101101100"),
								 ("1100001010110011","1110110110011100"),
								 ("1100001010100101","1110110111001100"),
								 ("1100001010010110","1110110111111100"),
								 ("1100001010001000","1110111000101101"),
								 ("1100001001111010","1110111001011101"),
								 ("1100001001101101","1110111010001101"),
								 ("1100001001011111","1110111010111110"),
								 ("1100001001010001","1110111011101110"),
								 ("1100001001000100","1110111100011111"),
								 ("1100001000110111","1110111101001111"),
								 ("1100001000101010","1110111110000000"),
								 ("1100001000011101","1110111110110000"),
								 ("1100001000010000","1110111111100001"),
								 ("1100001000000100","1111000000010010"),
								 ("1100000111110111","1111000001000010"),
								 ("1100000111101011","1111000001110011"),
								 ("1100000111011111","1111000010100100"),
								 ("1100000111010011","1111000011010101"),
								 ("1100000111000111","1111000100000101"),
								 ("1100000110111011","1111000100110110"),
								 ("1100000110110000","1111000101100111"),
								 ("1100000110100100","1111000110011000"),
								 ("1100000110011001","1111000111001001"),
								 ("1100000110001110","1111000111111010"),
								 ("1100000110000011","1111001000101011"),
								 ("1100000101111000","1111001001011100"),
								 ("1100000101101110","1111001010001110"),
								 ("1100000101100011","1111001010111111"),
								 ("1100000101011001","1111001011110000"),
								 ("1100000101001111","1111001100100001"),
								 ("1100000101000101","1111001101010010"),
								 ("1100000100111011","1111001110000100"),
								 ("1100000100110001","1111001110110101"),
								 ("1100000100101000","1111001111100110"),
								 ("1100000100011110","1111010000011000"),
								 ("1100000100010101","1111010001001001"),
								 ("1100000100001100","1111010001111011"),
								 ("1100000100000011","1111010010101100"),
								 ("1100000011111010","1111010011011101"),
								 ("1100000011110001","1111010100001111"),
								 ("1100000011101001","1111010101000000"),
								 ("1100000011100000","1111010101110010"),
								 ("1100000011011000","1111010110100100"),
								 ("1100000011010000","1111010111010101"),
								 ("1100000011001000","1111011000000111"),
								 ("1100000011000000","1111011000111001"),
								 ("1100000010111001","1111011001101010"),
								 ("1100000010110001","1111011010011100"),
								 ("1100000010101010","1111011011001110"),
								 ("1100000010100011","1111011011111111"),
								 ("1100000010011100","1111011100110001"),
								 ("1100000010010101","1111011101100011"),
								 ("1100000010001110","1111011110010101"),
								 ("1100000010001000","1111011111000111"),
								 ("1100000010000001","1111011111111001"),
								 ("1100000001111011","1111100000101010"),
								 ("1100000001110101","1111100001011100"),
								 ("1100000001101111","1111100010001110"),
								 ("1100000001101001","1111100011000000"),
								 ("1100000001100100","1111100011110010"),
								 ("1100000001011110","1111100100100100"),
								 ("1100000001011001","1111100101010110"),
								 ("1100000001010100","1111100110001000"),
								 ("1100000001001111","1111100110111010"),
								 ("1100000001001010","1111100111101100"),
								 ("1100000001000101","1111101000011110"),
								 ("1100000001000001","1111101001010000"),
								 ("1100000000111100","1111101010000010"),
								 ("1100000000111000","1111101010110100"),
								 ("1100000000110100","1111101011100110"),
								 ("1100000000110000","1111101100011001"),
								 ("1100000000101100","1111101101001011"),
								 ("1100000000101001","1111101101111101"),
								 ("1100000000100101","1111101110101111"),
								 ("1100000000100010","1111101111100001"),
								 ("1100000000011111","1111110000010011"),
								 ("1100000000011100","1111110001000101"),
								 ("1100000000011001","1111110001111000"),
								 ("1100000000010110","1111110010101010"),
								 ("1100000000010100","1111110011011100"),
								 ("1100000000010001","1111110100001110"),
								 ("1100000000001111","1111110101000000"),
								 ("1100000000001101","1111110101110011"),
								 ("1100000000001011","1111110110100101"),
								 ("1100000000001001","1111110111010111"),
								 ("1100000000001000","1111111000001001"),
								 ("1100000000000110","1111111000111100"),
								 ("1100000000000101","1111111001101110"),
								 ("1100000000000100","1111111010100000"),
								 ("1100000000000011","1111111011010010"),
								 ("1100000000000010","1111111100000101"),
								 ("1100000000000001","1111111100110111"),
								 ("1100000000000001","1111111101101001"),
								 ("1100000000000000","1111111110011011"),
								 ("1100000000000000","1111111111001110"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","1111111111100111"),
								 ("0100000000000000","1111111111001110"),
								 ("0100000000000000","1111111110110101"),
								 ("0100000000000000","1111111110011011"),
								 ("0100000000000000","1111111110000010"),
								 ("0011111111111111","1111111101101001"),
								 ("0011111111111111","1111111101010000"),
								 ("0011111111111111","1111111100110111"),
								 ("0011111111111110","1111111100011110"),
								 ("0011111111111110","1111111100000101"),
								 ("0011111111111110","1111111011101100"),
								 ("0011111111111101","1111111011010010"),
								 ("0011111111111101","1111111010111001"),
								 ("0011111111111100","1111111010100000"),
								 ("0011111111111100","1111111010000111"),
								 ("0011111111111011","1111111001101110"),
								 ("0011111111111010","1111111001010101"),
								 ("0011111111111010","1111111000111100"),
								 ("0011111111111001","1111111000100011"),
								 ("0011111111111000","1111111000001001"),
								 ("0011111111110111","1111110111110000"),
								 ("0011111111110111","1111110111010111"),
								 ("0011111111110110","1111110110111110"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111110100","1111110110001100"),
								 ("0011111111110011","1111110101110011"),
								 ("0011111111110010","1111110101011010"),
								 ("0011111111110001","1111110101000000"),
								 ("0011111111110000","1111110100100111"),
								 ("0011111111101111","1111110100001110"),
								 ("0011111111101101","1111110011110101"),
								 ("0011111111101100","1111110011011100"),
								 ("0011111111101011","1111110011000011"),
								 ("0011111111101010","1111110010101010"),
								 ("0011111111101000","1111110010010001"),
								 ("0011111111100111","1111110001111000"),
								 ("0011111111100110","1111110001011111"),
								 ("0011111111100100","1111110001000101"),
								 ("0011111111100011","1111110000101100"),
								 ("0011111111100001","1111110000010011"),
								 ("0011111111100000","1111101111111010"),
								 ("0011111111011110","1111101111100001"),
								 ("0011111111011100","1111101111001000"),
								 ("0011111111011011","1111101110101111"),
								 ("0011111111011001","1111101110010110"),
								 ("0011111111010111","1111101101111101"),
								 ("0011111111010101","1111101101100100"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111111010010","1111101100110010"),
								 ("0011111111010000","1111101100011001"),
								 ("0011111111001110","1111101100000000"),
								 ("0011111111001100","1111101011100110"),
								 ("0011111111001010","1111101011001101"),
								 ("0011111111001000","1111101010110100"),
								 ("0011111111000110","1111101010011011"),
								 ("0011111111000100","1111101010000010"),
								 ("0011111111000001","1111101001101001"),
								 ("0011111110111111","1111101001010000"),
								 ("0011111110111101","1111101000110111"),
								 ("0011111110111011","1111101000011110"),
								 ("0011111110111000","1111101000000101"),
								 ("0011111110110110","1111100111101100"),
								 ("0011111110110100","1111100111010011"),
								 ("0011111110110001","1111100110111010"),
								 ("0011111110101111","1111100110100001"),
								 ("0011111110101100","1111100110001000"),
								 ("0011111110101010","1111100101101111"),
								 ("0011111110100111","1111100101010110"),
								 ("0011111110100100","1111100100111101"),
								 ("0011111110100010","1111100100100100"),
								 ("0011111110011111","1111100100001011"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111110011001","1111100011011001"),
								 ("0011111110010111","1111100011000000"),
								 ("0011111110010100","1111100010100111"),
								 ("0011111110010001","1111100010001110"),
								 ("0011111110001110","1111100001110101"),
								 ("0011111110001011","1111100001011100"),
								 ("0011111110001000","1111100001000011"),
								 ("0011111110000101","1111100000101010"),
								 ("0011111110000010","1111100000010001"),
								 ("0011111101111111","1111011111111001"),
								 ("0011111101111011","1111011111100000"),
								 ("0011111101111000","1111011111000111"),
								 ("0011111101110101","1111011110101110"),
								 ("0011111101110010","1111011110010101"),
								 ("0011111101101110","1111011101111100"),
								 ("0011111101101011","1111011101100011"),
								 ("0011111101101000","1111011101001010"),
								 ("0011111101100100","1111011100110001"),
								 ("0011111101100001","1111011100011000"),
								 ("0011111101011101","1111011011111111"),
								 ("0011111101011010","1111011011100111"),
								 ("0011111101010110","1111011011001110"),
								 ("0011111101010010","1111011010110101"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111101001011","1111011010000011"),
								 ("0011111101000111","1111011001101010"),
								 ("0011111101000011","1111011001010001"),
								 ("0011111101000000","1111011000111001"),
								 ("0011111100111100","1111011000100000"),
								 ("0011111100111000","1111011000000111"),
								 ("0011111100110100","1111010111101110"),
								 ("0011111100110000","1111010111010101"),
								 ("0011111100101100","1111010110111100"),
								 ("0011111100101000","1111010110100100"),
								 ("0011111100100100","1111010110001011"),
								 ("0011111100100000","1111010101110010"),
								 ("0011111100011100","1111010101011001"),
								 ("0011111100010111","1111010101000000"),
								 ("0011111100010011","1111010100101000"),
								 ("0011111100001111","1111010100001111"),
								 ("0011111100001010","1111010011110110"),
								 ("0011111100000110","1111010011011101"),
								 ("0011111100000010","1111010011000101"),
								 ("0011111011111101","1111010010101100"),
								 ("0011111011111001","1111010010010011"),
								 ("0011111011110100","1111010001111011"),
								 ("0011111011110000","1111010001100010"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111011100111","1111010000110000"),
								 ("0011111011100010","1111010000011000"),
								 ("0011111011011101","1111001111111111"),
								 ("0011111011011000","1111001111100110"),
								 ("0011111011010100","1111001111001110"),
								 ("0011111011001111","1111001110110101"),
								 ("0011111011001010","1111001110011100"),
								 ("0011111011000101","1111001110000100"),
								 ("0011111011000000","1111001101101011"),
								 ("0011111010111011","1111001101010010"),
								 ("0011111010110110","1111001100111010"),
								 ("0011111010110001","1111001100100001"),
								 ("0011111010101100","1111001100001000"),
								 ("0011111010100111","1111001011110000"),
								 ("0011111010100010","1111001011010111"),
								 ("0011111010011101","1111001010111111"),
								 ("0011111010011000","1111001010100110"),
								 ("0011111010010010","1111001010001110"),
								 ("0011111010001101","1111001001110101"),
								 ("0011111010001000","1111001001011100"),
								 ("0011111010000010","1111001001000100"),
								 ("0011111001111101","1111001000101011"),
								 ("0011111001110111","1111001000010011"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111001101100","1111000111100010"),
								 ("0011111001100111","1111000111001001"),
								 ("0011111001100001","1111000110110001"),
								 ("0011111001011100","1111000110011000"),
								 ("0011111001010110","1111000110000000"),
								 ("0011111001010000","1111000101100111"),
								 ("0011111001001010","1111000101001111"),
								 ("0011111001000101","1111000100110110"),
								 ("0011111000111111","1111000100011110"),
								 ("0011111000111001","1111000100000101"),
								 ("0011111000110011","1111000011101101"),
								 ("0011111000101101","1111000011010101"),
								 ("0011111000100111","1111000010111100"),
								 ("0011111000100001","1111000010100100"),
								 ("0011111000011011","1111000010001011"),
								 ("0011111000010101","1111000001110011"),
								 ("0011111000001111","1111000001011011"),
								 ("0011111000001001","1111000001000010"),
								 ("0011111000000011","1111000000101010"),
								 ("0011110111111100","1111000000010010"),
								 ("0011110111110110","1110111111111001"),
								 ("0011110111110000","1110111111100001"),
								 ("0011110111101001","1110111111001001"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110111011101","1110111110011000"),
								 ("0011110111010110","1110111110000000"),
								 ("0011110111010000","1110111101100111"),
								 ("0011110111001001","1110111101001111"),
								 ("0011110111000010","1110111100110111"),
								 ("0011110110111100","1110111100011111"),
								 ("0011110110110101","1110111100000110"),
								 ("0011110110101111","1110111011101110"),
								 ("0011110110101000","1110111011010110"),
								 ("0011110110100001","1110111010111110"),
								 ("0011110110011010","1110111010100110"),
								 ("0011110110010011","1110111010001101"),
								 ("0011110110001101","1110111001110101"),
								 ("0011110110000110","1110111001011101"),
								 ("0011110101111111","1110111001000101"),
								 ("0011110101111000","1110111000101101"),
								 ("0011110101110001","1110111000010101"),
								 ("0011110101101010","1110110111111100"),
								 ("0011110101100011","1110110111100100"),
								 ("0011110101011011","1110110111001100"),
								 ("0011110101010100","1110110110110100"),
								 ("0011110101001101","1110110110011100"),
								 ("0011110101000110","1110110110000100"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110100110111","1110110101010100"),
								 ("0011110100110000","1110110100111100"),
								 ("0011110100101000","1110110100100100"),
								 ("0011110100100001","1110110100001100"),
								 ("0011110100011010","1110110011110100"),
								 ("0011110100010010","1110110011011100"),
								 ("0011110100001011","1110110011000100"),
								 ("0011110100000011","1110110010101100"),
								 ("0011110011111011","1110110010010100"),
								 ("0011110011110100","1110110001111100"),
								 ("0011110011101100","1110110001100100"),
								 ("0011110011100100","1110110001001100"),
								 ("0011110011011101","1110110000110100"),
								 ("0011110011010101","1110110000011100"),
								 ("0011110011001101","1110110000000101"),
								 ("0011110011000101","1110101111101101"),
								 ("0011110010111101","1110101111010101"),
								 ("0011110010110101","1110101110111101"),
								 ("0011110010101101","1110101110100101"),
								 ("0011110010100101","1110101110001101"),
								 ("0011110010011101","1110101101110101"),
								 ("0011110010010101","1110101101011110"),
								 ("0011110010001101","1110101101000110"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110001111101","1110101100010110"),
								 ("0011110001110100","1110101011111111"),
								 ("0011110001101100","1110101011100111"),
								 ("0011110001100100","1110101011001111"),
								 ("0011110001011011","1110101010110111"),
								 ("0011110001010011","1110101010100000"),
								 ("0011110001001011","1110101010001000"),
								 ("0011110001000010","1110101001110000"),
								 ("0011110000111010","1110101001011001"),
								 ("0011110000110001","1110101001000001"),
								 ("0011110000101001","1110101000101001"),
								 ("0011110000100000","1110101000010010"),
								 ("0011110000010111","1110100111111010"),
								 ("0011110000001111","1110100111100011"),
								 ("0011110000000110","1110100111001011"),
								 ("0011101111111101","1110100110110100"),
								 ("0011101111110101","1110100110011100"),
								 ("0011101111101100","1110100110000100"),
								 ("0011101111100011","1110100101101101"),
								 ("0011101111011010","1110100101010101"),
								 ("0011101111010001","1110100100111110"),
								 ("0011101111001000","1110100100100110"),
								 ("0011101110111111","1110100100001111"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101110101101","1110100011100000"),
								 ("0011101110100100","1110100011001001"),
								 ("0011101110011011","1110100010110001"),
								 ("0011101110010010","1110100010011010"),
								 ("0011101110001000","1110100010000010"),
								 ("0011101101111111","1110100001101011"),
								 ("0011101101110110","1110100001010100"),
								 ("0011101101101101","1110100000111100"),
								 ("0011101101100011","1110100000100101"),
								 ("0011101101011010","1110100000001110"),
								 ("0011101101010000","1110011111110110"),
								 ("0011101101000111","1110011111011111"),
								 ("0011101100111110","1110011111001000"),
								 ("0011101100110100","1110011110110001"),
								 ("0011101100101010","1110011110011001"),
								 ("0011101100100001","1110011110000010"),
								 ("0011101100010111","1110011101101011"),
								 ("0011101100001110","1110011101010100"),
								 ("0011101100000100","1110011100111101"),
								 ("0011101011111010","1110011100100101"),
								 ("0011101011110000","1110011100001110"),
								 ("0011101011100110","1110011011110111"),
								 ("0011101011011101","1110011011100000"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101011001001","1110011010110010"),
								 ("0011101010111111","1110011010011011"),
								 ("0011101010110101","1110011010000100"),
								 ("0011101010101011","1110011001101101"),
								 ("0011101010100001","1110011001010110"),
								 ("0011101010010111","1110011000111111"),
								 ("0011101010001101","1110011000101000"),
								 ("0011101010000010","1110011000010001"),
								 ("0011101001111000","1110010111111010"),
								 ("0011101001101110","1110010111100011"),
								 ("0011101001100100","1110010111001100"),
								 ("0011101001011001","1110010110110101"),
								 ("0011101001001111","1110010110011110"),
								 ("0011101001000101","1110010110000111"),
								 ("0011101000111010","1110010101110000"),
								 ("0011101000110000","1110010101011001"),
								 ("0011101000100101","1110010101000010"),
								 ("0011101000011011","1110010100101100"),
								 ("0011101000010000","1110010100010101"),
								 ("0011101000000110","1110010011111110"),
								 ("0011100111111011","1110010011100111"),
								 ("0011100111110000","1110010011010000"),
								 ("0011100111100110","1110010010111010"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100111010000","1110010010001100"),
								 ("0011100111000101","1110010001110110"),
								 ("0011100110111011","1110010001011111"),
								 ("0011100110110000","1110010001001000"),
								 ("0011100110100101","1110010000110010"),
								 ("0011100110011010","1110010000011011"),
								 ("0011100110001111","1110010000000100"),
								 ("0011100110000100","1110001111101110"),
								 ("0011100101111001","1110001111010111"),
								 ("0011100101101110","1110001111000001"),
								 ("0011100101100011","1110001110101010"),
								 ("0011100101011000","1110001110010100"),
								 ("0011100101001100","1110001101111101"),
								 ("0011100101000001","1110001101100111"),
								 ("0011100100110110","1110001101010000"),
								 ("0011100100101011","1110001100111010"),
								 ("0011100100011111","1110001100100011"),
								 ("0011100100010100","1110001100001101"),
								 ("0011100100001001","1110001011110110"),
								 ("0011100011111101","1110001011100000"),
								 ("0011100011110010","1110001011001010"),
								 ("0011100011100110","1110001010110011"),
								 ("0011100011011011","1110001010011101"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100011000011","1110001001110000"),
								 ("0011100010111000","1110001001011010"),
								 ("0011100010101100","1110001001000100"),
								 ("0011100010100001","1110001000101101"),
								 ("0011100010010101","1110001000010111"),
								 ("0011100010001001","1110001000000001"),
								 ("0011100001111101","1110000111101011"),
								 ("0011100001110001","1110000111010101"),
								 ("0011100001100110","1110000110111110"),
								 ("0011100001011010","1110000110101000"),
								 ("0011100001001110","1110000110010010"),
								 ("0011100001000010","1110000101111100"),
								 ("0011100000110110","1110000101100110"),
								 ("0011100000101010","1110000101010000"),
								 ("0011100000011110","1110000100111010"),
								 ("0011100000010010","1110000100100100"),
								 ("0011100000000101","1110000100001110"),
								 ("0011011111111001","1110000011111000"),
								 ("0011011111101101","1110000011100010"),
								 ("0011011111100001","1110000011001100"),
								 ("0011011111010101","1110000010110110"),
								 ("0011011111001000","1110000010100000"),
								 ("0011011110111100","1110000010001010"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011110100011","1110000001011110"),
								 ("0011011110010111","1110000001001001"),
								 ("0011011110001010","1110000000110011"),
								 ("0011011101111110","1110000000011101"),
								 ("0011011101110001","1110000000000111"),
								 ("0011011101100101","1101111111110001"),
								 ("0011011101011000","1101111111011100"),
								 ("0011011101001011","1101111111000110"),
								 ("0011011100111111","1101111110110000"),
								 ("0011011100110010","1101111110011011"),
								 ("0011011100100101","1101111110000101"),
								 ("0011011100011000","1101111101101111"),
								 ("0011011100001100","1101111101011010"),
								 ("0011011011111111","1101111101000100"),
								 ("0011011011110010","1101111100101111"),
								 ("0011011011100101","1101111100011001"),
								 ("0011011011011000","1101111100000011"),
								 ("0011011011001011","1101111011101110"),
								 ("0011011010111110","1101111011011000"),
								 ("0011011010110001","1101111011000011"),
								 ("0011011010100100","1101111010101101"),
								 ("0011011010010111","1101111010011000"),
								 ("0011011010001010","1101111010000011"),
								 ("0011011001111101","1101111001101101"),
								 ("0011011001101111","1101111001011000"),
								 ("0011011001100010","1101111001000010"),
								 ("0011011001010101","1101111000101101"),
								 ("0011011001001000","1101111000011000"),
								 ("0011011000111010","1101111000000010"),
								 ("0011011000101101","1101110111101101"),
								 ("0011011000100000","1101110111011000"),
								 ("0011011000010010","1101110111000011"),
								 ("0011011000000101","1101110110101101"),
								 ("0011010111110111","1101110110011000"),
								 ("0011010111101010","1101110110000011"),
								 ("0011010111011100","1101110101101110"),
								 ("0011010111001110","1101110101011001"),
								 ("0011010111000001","1101110101000100"),
								 ("0011010110110011","1101110100101110"),
								 ("0011010110100101","1101110100011001"),
								 ("0011010110011000","1101110100000100"),
								 ("0011010110001010","1101110011101111"),
								 ("0011010101111100","1101110011011010"),
								 ("0011010101101110","1101110011000101"),
								 ("0011010101100001","1101110010110000"),
								 ("0011010101010011","1101110010011011"),
								 ("0011010101000101","1101110010000110"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010100101001","1101110001011101"),
								 ("0011010100011011","1101110001001000"),
								 ("0011010100001101","1101110000110011"),
								 ("0011010011111111","1101110000011110"),
								 ("0011010011110001","1101110000001001"),
								 ("0011010011100010","1101101111110101"),
								 ("0011010011010100","1101101111100000"),
								 ("0011010011000110","1101101111001011"),
								 ("0011010010111000","1101101110110110"),
								 ("0011010010101010","1101101110100010"),
								 ("0011010010011011","1101101110001101"),
								 ("0011010010001101","1101101101111000"),
								 ("0011010001111111","1101101101100100"),
								 ("0011010001110000","1101101101001111"),
								 ("0011010001100010","1101101100111011"),
								 ("0011010001010011","1101101100100110"),
								 ("0011010001000101","1101101100010001"),
								 ("0011010000110110","1101101011111101"),
								 ("0011010000101000","1101101011101000"),
								 ("0011010000011001","1101101011010100"),
								 ("0011010000001011","1101101010111111"),
								 ("0011001111111100","1101101010101011"),
								 ("0011001111101101","1101101010010111"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001111010000","1101101001101110"),
								 ("0011001111000001","1101101001011010"),
								 ("0011001110110010","1101101001000101"),
								 ("0011001110100011","1101101000110001"),
								 ("0011001110010101","1101101000011101"),
								 ("0011001110000110","1101101000001000"),
								 ("0011001101110111","1101100111110100"),
								 ("0011001101101000","1101100111100000"),
								 ("0011001101011001","1101100111001100"),
								 ("0011001101001010","1101100110111000"),
								 ("0011001100111011","1101100110100100"),
								 ("0011001100101100","1101100110001111"),
								 ("0011001100011101","1101100101111011"),
								 ("0011001100001101","1101100101100111"),
								 ("0011001011111110","1101100101010011"),
								 ("0011001011101111","1101100100111111"),
								 ("0011001011100000","1101100100101011"),
								 ("0011001011010000","1101100100010111"),
								 ("0011001011000001","1101100100000011"),
								 ("0011001010110010","1101100011101111"),
								 ("0011001010100011","1101100011011100"),
								 ("0011001010010011","1101100011001000"),
								 ("0011001010000100","1101100010110100"),
								 ("0011001001110100","1101100010100000"),
								 ("0011001001100101","1101100010001100"),
								 ("0011001001010101","1101100001111000"),
								 ("0011001001000110","1101100001100101"),
								 ("0011001000110110","1101100001010001"),
								 ("0011001000100111","1101100000111101"),
								 ("0011001000010111","1101100000101010"),
								 ("0011001000000111","1101100000010110"),
								 ("0011000111111000","1101100000000010"),
								 ("0011000111101000","1101011111101111"),
								 ("0011000111011000","1101011111011011"),
								 ("0011000111001000","1101011111001000"),
								 ("0011000110111001","1101011110110100"),
								 ("0011000110101001","1101011110100000"),
								 ("0011000110011001","1101011110001101"),
								 ("0011000110001001","1101011101111010"),
								 ("0011000101111001","1101011101100110"),
								 ("0011000101101001","1101011101010011"),
								 ("0011000101011001","1101011100111111"),
								 ("0011000101001001","1101011100101100"),
								 ("0011000100111001","1101011100011001"),
								 ("0011000100101001","1101011100000101"),
								 ("0011000100011001","1101011011110010"),
								 ("0011000100001001","1101011011011111"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000011101000","1101011010111000"),
								 ("0011000011011000","1101011010100101"),
								 ("0011000011001000","1101011010010010"),
								 ("0011000010111000","1101011001111111"),
								 ("0011000010100111","1101011001101100"),
								 ("0011000010010111","1101011001011001"),
								 ("0011000010000111","1101011001000101"),
								 ("0011000001110110","1101011000110010"),
								 ("0011000001100110","1101011000011111"),
								 ("0011000001010101","1101011000001100"),
								 ("0011000001000101","1101010111111001"),
								 ("0011000000110100","1101010111100110"),
								 ("0011000000100100","1101010111010100"),
								 ("0011000000010011","1101010111000001"),
								 ("0011000000000010","1101010110101110"),
								 ("0010111111110010","1101010110011011"),
								 ("0010111111100001","1101010110001000"),
								 ("0010111111010000","1101010101110101"),
								 ("0010111111000000","1101010101100011"),
								 ("0010111110101111","1101010101010000"),
								 ("0010111110011110","1101010100111101"),
								 ("0010111110001101","1101010100101010"),
								 ("0010111101111101","1101010100011000"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111101011011","1101010011110011"),
								 ("0010111101001010","1101010011100000"),
								 ("0010111100111001","1101010011001101"),
								 ("0010111100101000","1101010010111011"),
								 ("0010111100010111","1101010010101000"),
								 ("0010111100000110","1101010010010110"),
								 ("0010111011110101","1101010010000011"),
								 ("0010111011100100","1101010001110001"),
								 ("0010111011010011","1101010001011111"),
								 ("0010111011000010","1101010001001100"),
								 ("0010111010110000","1101010000111010"),
								 ("0010111010011111","1101010000101000"),
								 ("0010111010001110","1101010000010101"),
								 ("0010111001111101","1101010000000011"),
								 ("0010111001101011","1101001111110001"),
								 ("0010111001011010","1101001111011111"),
								 ("0010111001001001","1101001111001100"),
								 ("0010111000110111","1101001110111010"),
								 ("0010111000100110","1101001110101000"),
								 ("0010111000010101","1101001110010110"),
								 ("0010111000000011","1101001110000100"),
								 ("0010110111110010","1101001101110010"),
								 ("0010110111100000","1101001101100000"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110110111101","1101001100111100"),
								 ("0010110110101011","1101001100101010"),
								 ("0010110110011010","1101001100011000"),
								 ("0010110110001000","1101001100000110"),
								 ("0010110101110110","1101001011110100"),
								 ("0010110101100101","1101001011100010"),
								 ("0010110101010011","1101001011010001"),
								 ("0010110101000001","1101001010111111"),
								 ("0010110100101111","1101001010101101"),
								 ("0010110100011110","1101001010011011"),
								 ("0010110100001100","1101001010001010"),
								 ("0010110011111010","1101001001111000"),
								 ("0010110011101000","1101001001100110"),
								 ("0010110011010110","1101001001010101"),
								 ("0010110011000100","1101001001000011"),
								 ("0010110010110010","1101001000110001"),
								 ("0010110010100000","1101001000100000"),
								 ("0010110010001110","1101001000001110"),
								 ("0010110001111100","1101000111111101"),
								 ("0010110001101010","1101000111101011"),
								 ("0010110001011000","1101000111011010"),
								 ("0010110001000110","1101000111001001"),
								 ("0010110000110100","1101000110110111"),
								 ("0010110000100001","1101000110100110"),
								 ("0010110000001111","1101000110010101"),
								 ("0010101111111101","1101000110000011"),
								 ("0010101111101011","1101000101110010"),
								 ("0010101111011000","1101000101100001"),
								 ("0010101111000110","1101000101010000"),
								 ("0010101110110100","1101000100111110"),
								 ("0010101110100001","1101000100101101"),
								 ("0010101110001111","1101000100011100"),
								 ("0010101101111101","1101000100001011"),
								 ("0010101101101010","1101000011111010"),
								 ("0010101101011000","1101000011101001"),
								 ("0010101101000101","1101000011011000"),
								 ("0010101100110011","1101000011000111"),
								 ("0010101100100000","1101000010110110"),
								 ("0010101100001101","1101000010100101"),
								 ("0010101011111011","1101000010010100"),
								 ("0010101011101000","1101000010000011"),
								 ("0010101011010110","1101000001110011"),
								 ("0010101011000011","1101000001100010"),
								 ("0010101010110000","1101000001010001"),
								 ("0010101010011101","1101000001000000"),
								 ("0010101010001011","1101000000110000"),
								 ("0010101001111000","1101000000011111"),
								 ("0010101001100101","1101000000001110"),
								 ("0010101001010010","1100111111111110"),
								 ("0010101000111111","1100111111101101"),
								 ("0010101000101100","1100111111011100"),
								 ("0010101000011010","1100111111001100"),
								 ("0010101000000111","1100111110111011"),
								 ("0010100111110100","1100111110101011"),
								 ("0010100111100001","1100111110011010"),
								 ("0010100111001110","1100111110001010"),
								 ("0010100110111011","1100111101111001"),
								 ("0010100110100111","1100111101101001"),
								 ("0010100110010100","1100111101011001"),
								 ("0010100110000001","1100111101001000"),
								 ("0010100101101110","1100111100111000"),
								 ("0010100101011011","1100111100101000"),
								 ("0010100101001000","1100111100011000"),
								 ("0010100100110101","1100111100000111"),
								 ("0010100100100001","1100111011110111"),
								 ("0010100100001110","1100111011100111"),
								 ("0010100011111011","1100111011010111"),
								 ("0010100011100111","1100111011000111"),
								 ("0010100011010100","1100111010110111"),
								 ("0010100011000001","1100111010100111"),
								 ("0010100010101101","1100111010010111"),
								 ("0010100010011010","1100111010000111"),
								 ("0010100010000110","1100111001110111"),
								 ("0010100001110011","1100111001100111"),
								 ("0010100001100000","1100111001010111"),
								 ("0010100001001100","1100111001000111"),
								 ("0010100000111000","1100111000111000"),
								 ("0010100000100101","1100111000101000"),
								 ("0010100000010001","1100111000011000"),
								 ("0010011111111110","1100111000001000"),
								 ("0010011111101010","1100110111111001"),
								 ("0010011111010110","1100110111101001"),
								 ("0010011111000011","1100110111011001"),
								 ("0010011110101111","1100110111001010"),
								 ("0010011110011011","1100110110111010"),
								 ("0010011110001000","1100110110101011"),
								 ("0010011101110100","1100110110011011"),
								 ("0010011101100000","1100110110001100"),
								 ("0010011101001100","1100110101111100"),
								 ("0010011100111000","1100110101101101"),
								 ("0010011100100100","1100110101011101"),
								 ("0010011100010001","1100110101001110"),
								 ("0010011011111101","1100110100111111"),
								 ("0010011011101001","1100110100110000"),
								 ("0010011011010101","1100110100100000"),
								 ("0010011011000001","1100110100010001"),
								 ("0010011010101101","1100110100000010"),
								 ("0010011010011001","1100110011110011"),
								 ("0010011010000101","1100110011100011"),
								 ("0010011001110001","1100110011010100"),
								 ("0010011001011100","1100110011000101"),
								 ("0010011001001000","1100110010110110"),
								 ("0010011000110100","1100110010100111"),
								 ("0010011000100000","1100110010011000"),
								 ("0010011000001100","1100110010001001"),
								 ("0010010111111000","1100110001111010"),
								 ("0010010111100011","1100110001101011"),
								 ("0010010111001111","1100110001011101"),
								 ("0010010110111011","1100110001001110"),
								 ("0010010110100110","1100110000111111"),
								 ("0010010110010010","1100110000110000"),
								 ("0010010101111110","1100110000100001"),
								 ("0010010101101001","1100110000010011"),
								 ("0010010101010101","1100110000000100"),
								 ("0010010101000001","1100101111110101"),
								 ("0010010100101100","1100101111100111"),
								 ("0010010100011000","1100101111011000"),
								 ("0010010100000011","1100101111001010"),
								 ("0010010011101111","1100101110111011"),
								 ("0010010011011010","1100101110101101"),
								 ("0010010011000101","1100101110011110"),
								 ("0010010010110001","1100101110010000"),
								 ("0010010010011100","1100101110000001"),
								 ("0010010010001000","1100101101110011"),
								 ("0010010001110011","1100101101100101"),
								 ("0010010001011110","1100101101010110"),
								 ("0010010001001010","1100101101001000"),
								 ("0010010000110101","1100101100111010"),
								 ("0010010000100000","1100101100101100"),
								 ("0010010000001011","1100101100011110"),
								 ("0010001111110111","1100101100001111"),
								 ("0010001111100010","1100101100000001"),
								 ("0010001111001101","1100101011110011"),
								 ("0010001110111000","1100101011100101"),
								 ("0010001110100011","1100101011010111"),
								 ("0010001110001110","1100101011001001"),
								 ("0010001101111010","1100101010111011"),
								 ("0010001101100101","1100101010101101"),
								 ("0010001101010000","1100101010011111"),
								 ("0010001100111011","1100101010010010"),
								 ("0010001100100110","1100101010000100"),
								 ("0010001100010001","1100101001110110"),
								 ("0010001011111100","1100101001101000"),
								 ("0010001011100111","1100101001011011"),
								 ("0010001011010010","1100101001001101"),
								 ("0010001010111100","1100101000111111"),
								 ("0010001010100111","1100101000110010"),
								 ("0010001010010010","1100101000100100"),
								 ("0010001001111101","1100101000010110"),
								 ("0010001001101000","1100101000001001"),
								 ("0010001001010011","1100100111111011"),
								 ("0010001000111101","1100100111101110"),
								 ("0010001000101000","1100100111100000"),
								 ("0010001000010011","1100100111010011"),
								 ("0010000111111110","1100100111000110"),
								 ("0010000111101000","1100100110111000"),
								 ("0010000111010011","1100100110101011"),
								 ("0010000110111110","1100100110011110"),
								 ("0010000110101000","1100100110010001"),
								 ("0010000110010011","1100100110000011"),
								 ("0010000101111101","1100100101110110"),
								 ("0010000101101000","1100100101101001"),
								 ("0010000101010011","1100100101011100"),
								 ("0010000100111101","1100100101001111"),
								 ("0010000100101000","1100100101000010"),
								 ("0010000100010010","1100100100110101"),
								 ("0010000011111101","1100100100101000"),
								 ("0010000011100111","1100100100011011"),
								 ("0010000011010001","1100100100001110"),
								 ("0010000010111100","1100100100000001"),
								 ("0010000010100110","1100100011110100"),
								 ("0010000010010001","1100100011101000"),
								 ("0010000001111011","1100100011011011"),
								 ("0010000001100101","1100100011001110"),
								 ("0010000001010000","1100100011000001"),
								 ("0010000000111010","1100100010110101"),
								 ("0010000000100100","1100100010101000"),
								 ("0010000000001111","1100100010011011"),
								 ("0001111111111001","1100100010001111"),
								 ("0001111111100011","1100100010000010"),
								 ("0001111111001101","1100100001110110"),
								 ("0001111110110111","1100100001101001"),
								 ("0001111110100010","1100100001011101"),
								 ("0001111110001100","1100100001010000"),
								 ("0001111101110110","1100100001000100"),
								 ("0001111101100000","1100100000111000"),
								 ("0001111101001010","1100100000101011"),
								 ("0001111100110100","1100100000011111"),
								 ("0001111100011110","1100100000010011"),
								 ("0001111100001000","1100100000000111"),
								 ("0001111011110010","1100011111111011"),
								 ("0001111011011100","1100011111101110"),
								 ("0001111011000110","1100011111100010"),
								 ("0001111010110000","1100011111010110"),
								 ("0001111010011010","1100011111001010"),
								 ("0001111010000100","1100011110111110"),
								 ("0001111001101110","1100011110110010"),
								 ("0001111001011000","1100011110100110"),
								 ("0001111001000010","1100011110011010"),
								 ("0001111000101011","1100011110001111"),
								 ("0001111000010101","1100011110000011"),
								 ("0001110111111111","1100011101110111"),
								 ("0001110111101001","1100011101101011"),
								 ("0001110111010011","1100011101011111"),
								 ("0001110110111100","1100011101010100"),
								 ("0001110110100110","1100011101001000"),
								 ("0001110110010000","1100011100111101"),
								 ("0001110101111001","1100011100110001"),
								 ("0001110101100011","1100011100100101"),
								 ("0001110101001101","1100011100011010"),
								 ("0001110100110110","1100011100001110"),
								 ("0001110100100000","1100011100000011"),
								 ("0001110100001010","1100011011110111"),
								 ("0001110011110011","1100011011101100"),
								 ("0001110011011101","1100011011100001"),
								 ("0001110011000110","1100011011010101"),
								 ("0001110010110000","1100011011001010"),
								 ("0001110010011001","1100011010111111"),
								 ("0001110010000011","1100011010110100"),
								 ("0001110001101100","1100011010101000"),
								 ("0001110001010110","1100011010011101"),
								 ("0001110000111111","1100011010010010"),
								 ("0001110000101001","1100011010000111"),
								 ("0001110000010010","1100011001111100"),
								 ("0001101111111100","1100011001110001"),
								 ("0001101111100101","1100011001100110"),
								 ("0001101111001110","1100011001011011"),
								 ("0001101110111000","1100011001010000"),
								 ("0001101110100001","1100011001000101"),
								 ("0001101110001010","1100011000111011"),
								 ("0001101101110100","1100011000110000"),
								 ("0001101101011101","1100011000100101"),
								 ("0001101101000110","1100011000011010"),
								 ("0001101100110000","1100011000010000"),
								 ("0001101100011001","1100011000000101"),
								 ("0001101100000010","1100010111111010"),
								 ("0001101011101011","1100010111110000"),
								 ("0001101011010100","1100010111100101"),
								 ("0001101010111110","1100010111011011"),
								 ("0001101010100111","1100010111010000"),
								 ("0001101010010000","1100010111000110"),
								 ("0001101001111001","1100010110111011"),
								 ("0001101001100010","1100010110110001"),
								 ("0001101001001011","1100010110100111"),
								 ("0001101000110100","1100010110011100"),
								 ("0001101000011101","1100010110010010"),
								 ("0001101000000110","1100010110001000"),
								 ("0001100111101111","1100010101111110"),
								 ("0001100111011000","1100010101110011"),
								 ("0001100111000001","1100010101101001"),
								 ("0001100110101010","1100010101011111"),
								 ("0001100110010011","1100010101010101"),
								 ("0001100101111100","1100010101001011"),
								 ("0001100101100101","1100010101000001"),
								 ("0001100101001110","1100010100110111"),
								 ("0001100100110111","1100010100101101"),
								 ("0001100100100000","1100010100100011"),
								 ("0001100100001001","1100010100011010"),
								 ("0001100011110010","1100010100010000"),
								 ("0001100011011011","1100010100000110"),
								 ("0001100011000011","1100010011111100"),
								 ("0001100010101100","1100010011110010"),
								 ("0001100010010101","1100010011101001"),
								 ("0001100001111110","1100010011011111"),
								 ("0001100001100111","1100010011010110"),
								 ("0001100001001111","1100010011001100"),
								 ("0001100000111000","1100010011000010"),
								 ("0001100000100001","1100010010111001"),
								 ("0001100000001010","1100010010110000"),
								 ("0001011111110010","1100010010100110"),
								 ("0001011111011011","1100010010011101"),
								 ("0001011111000100","1100010010010011"),
								 ("0001011110101100","1100010010001010"),
								 ("0001011110010101","1100010010000001"),
								 ("0001011101111110","1100010001111000"),
								 ("0001011101100110","1100010001101110"),
								 ("0001011101001111","1100010001100101"),
								 ("0001011100110111","1100010001011100"),
								 ("0001011100100000","1100010001010011"),
								 ("0001011100001001","1100010001001010"),
								 ("0001011011110001","1100010001000001"),
								 ("0001011011011010","1100010000111000"),
								 ("0001011011000010","1100010000101111"),
								 ("0001011010101011","1100010000100110"),
								 ("0001011010010011","1100010000011101"),
								 ("0001011001111100","1100010000010100"),
								 ("0001011001100100","1100010000001011"),
								 ("0001011001001100","1100010000000011"),
								 ("0001011000110101","1100001111111010"),
								 ("0001011000011101","1100001111110001"),
								 ("0001011000000110","1100001111101001"),
								 ("0001010111101110","1100001111100000"),
								 ("0001010111010111","1100001111010111"),
								 ("0001010110111111","1100001111001111"),
								 ("0001010110100111","1100001111000110"),
								 ("0001010110010000","1100001110111110"),
								 ("0001010101111000","1100001110110101"),
								 ("0001010101100000","1100001110101101"),
								 ("0001010101001001","1100001110100101"),
								 ("0001010100110001","1100001110011100"),
								 ("0001010100011001","1100001110010100"),
								 ("0001010100000001","1100001110001100"),
								 ("0001010011101010","1100001110000011"),
								 ("0001010011010010","1100001101111011"),
								 ("0001010010111010","1100001101110011"),
								 ("0001010010100010","1100001101101011"),
								 ("0001010010001011","1100001101100011"),
								 ("0001010001110011","1100001101011011"),
								 ("0001010001011011","1100001101010011"),
								 ("0001010001000011","1100001101001011"),
								 ("0001010000101011","1100001101000011"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001111111011","1100001100110011"),
								 ("0001001111100100","1100001100101011"),
								 ("0001001111001100","1100001100100011"),
								 ("0001001110110100","1100001100011100"),
								 ("0001001110011100","1100001100010100"),
								 ("0001001110000100","1100001100001100"),
								 ("0001001101101100","1100001100000101"),
								 ("0001001101010100","1100001011111101"),
								 ("0001001100111100","1100001011110101"),
								 ("0001001100100100","1100001011101110"),
								 ("0001001100001100","1100001011100110"),
								 ("0001001011110100","1100001011011111"),
								 ("0001001011011100","1100001011011000"),
								 ("0001001011000100","1100001011010000"),
								 ("0001001010101100","1100001011001001"),
								 ("0001001010010100","1100001011000001"),
								 ("0001001001111100","1100001010111010"),
								 ("0001001001100100","1100001010110011"),
								 ("0001001001001100","1100001010101100"),
								 ("0001001000110100","1100001010100101"),
								 ("0001001000011100","1100001010011101"),
								 ("0001001000000100","1100001010010110"),
								 ("0001000111101011","1100001010001111"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000110111011","1100001010000001"),
								 ("0001000110100011","1100001001111010"),
								 ("0001000110001011","1100001001110011"),
								 ("0001000101110011","1100001001101101"),
								 ("0001000101011010","1100001001100110"),
								 ("0001000101000010","1100001001011111"),
								 ("0001000100101010","1100001001011000"),
								 ("0001000100010010","1100001001010001"),
								 ("0001000011111010","1100001001001011"),
								 ("0001000011100001","1100001001000100"),
								 ("0001000011001001","1100001000111110"),
								 ("0001000010110001","1100001000110111"),
								 ("0001000010011001","1100001000110000"),
								 ("0001000010000000","1100001000101010"),
								 ("0001000001101000","1100001000100011"),
								 ("0001000001010000","1100001000011101"),
								 ("0001000000110111","1100001000010111"),
								 ("0001000000011111","1100001000010000"),
								 ("0001000000000111","1100001000001010"),
								 ("0000111111101110","1100001000000100"),
								 ("0000111111010110","1100000111111101"),
								 ("0000111110111110","1100000111110111"),
								 ("0000111110100101","1100000111110001"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111101110101","1100000111100101"),
								 ("0000111101011100","1100000111011111"),
								 ("0000111101000100","1100000111011001"),
								 ("0000111100101011","1100000111010011"),
								 ("0000111100010011","1100000111001101"),
								 ("0000111011111011","1100000111000111"),
								 ("0000111011100010","1100000111000001"),
								 ("0000111011001010","1100000110111011"),
								 ("0000111010110001","1100000110110110"),
								 ("0000111010011001","1100000110110000"),
								 ("0000111010000000","1100000110101010"),
								 ("0000111001101000","1100000110100100"),
								 ("0000111001001111","1100000110011111"),
								 ("0000111000110111","1100000110011001"),
								 ("0000111000011110","1100000110010100"),
								 ("0000111000000110","1100000110001110"),
								 ("0000110111101101","1100000110001001"),
								 ("0000110111010101","1100000110000011"),
								 ("0000110110111100","1100000101111110"),
								 ("0000110110100100","1100000101111000"),
								 ("0000110110001011","1100000101110011"),
								 ("0000110101110010","1100000101101110"),
								 ("0000110101011010","1100000101101000"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110100101001","1100000101011110"),
								 ("0000110100010000","1100000101011001"),
								 ("0000110011111000","1100000101010100"),
								 ("0000110011011111","1100000101001111"),
								 ("0000110011000110","1100000101001010"),
								 ("0000110010101110","1100000101000101"),
								 ("0000110010010101","1100000101000000"),
								 ("0000110001111100","1100000100111011"),
								 ("0000110001100100","1100000100110110"),
								 ("0000110001001011","1100000100110001"),
								 ("0000110000110010","1100000100101100"),
								 ("0000110000011010","1100000100101000"),
								 ("0000110000000001","1100000100100011"),
								 ("0000101111101000","1100000100011110"),
								 ("0000101111010000","1100000100011001"),
								 ("0000101110110111","1100000100010101"),
								 ("0000101110011110","1100000100010000"),
								 ("0000101110000101","1100000100001100"),
								 ("0000101101101101","1100000100000111"),
								 ("0000101101010100","1100000100000011"),
								 ("0000101100111011","1100000011111110"),
								 ("0000101100100011","1100000011111010"),
								 ("0000101100001010","1100000011110110"),
								 ("0000101011110001","1100000011110001"),
								 ("0000101011011000","1100000011101101"),
								 ("0000101011000000","1100000011101001"),
								 ("0000101010100111","1100000011100100"),
								 ("0000101010001110","1100000011100000"),
								 ("0000101001110101","1100000011011100"),
								 ("0000101001011100","1100000011011000"),
								 ("0000101001000100","1100000011010100"),
								 ("0000101000101011","1100000011010000"),
								 ("0000101000010010","1100000011001100"),
								 ("0000100111111001","1100000011001000"),
								 ("0000100111100000","1100000011000100"),
								 ("0000100111000111","1100000011000000"),
								 ("0000100110101111","1100000010111101"),
								 ("0000100110010110","1100000010111001"),
								 ("0000100101111101","1100000010110101"),
								 ("0000100101100100","1100000010110001"),
								 ("0000100101001011","1100000010101110"),
								 ("0000100100110010","1100000010101010"),
								 ("0000100100011001","1100000010100110"),
								 ("0000100100000001","1100000010100011"),
								 ("0000100011101000","1100000010011111"),
								 ("0000100011001111","1100000010011100"),
								 ("0000100010110110","1100000010011000"),
								 ("0000100010011101","1100000010010101"),
								 ("0000100010000100","1100000010010010"),
								 ("0000100001101011","1100000010001110"),
								 ("0000100001010010","1100000010001011"),
								 ("0000100000111001","1100000010001000"),
								 ("0000100000100000","1100000010000101"),
								 ("0000100000000111","1100000010000001"),
								 ("0000011111101111","1100000001111110"),
								 ("0000011111010110","1100000001111011"),
								 ("0000011110111101","1100000001111000"),
								 ("0000011110100100","1100000001110101"),
								 ("0000011110001011","1100000001110010"),
								 ("0000011101110010","1100000001101111"),
								 ("0000011101011001","1100000001101100"),
								 ("0000011101000000","1100000001101001"),
								 ("0000011100100111","1100000001100111"),
								 ("0000011100001110","1100000001100100"),
								 ("0000011011110101","1100000001100001"),
								 ("0000011011011100","1100000001011110"),
								 ("0000011011000011","1100000001011100"),
								 ("0000011010101010","1100000001011001"),
								 ("0000011010010001","1100000001010110"),
								 ("0000011001111000","1100000001010100"),
								 ("0000011001011111","1100000001010001"),
								 ("0000011001000110","1100000001001111"),
								 ("0000011000101101","1100000001001100"),
								 ("0000011000010100","1100000001001010"),
								 ("0000010111111011","1100000001001000"),
								 ("0000010111100010","1100000001000101"),
								 ("0000010111001001","1100000001000011"),
								 ("0000010110110000","1100000001000001"),
								 ("0000010110010111","1100000000111111"),
								 ("0000010101111110","1100000000111100"),
								 ("0000010101100101","1100000000111010"),
								 ("0000010101001100","1100000000111000"),
								 ("0000010100110011","1100000000110110"),
								 ("0000010100011010","1100000000110100"),
								 ("0000010100000000","1100000000110010"),
								 ("0000010011100111","1100000000110000"),
								 ("0000010011001110","1100000000101110"),
								 ("0000010010110101","1100000000101100"),
								 ("0000010010011100","1100000000101011"),
								 ("0000010010000011","1100000000101001"),
								 ("0000010001101010","1100000000100111"),
								 ("0000010001010001","1100000000100101"),
								 ("0000010000111000","1100000000100100"),
								 ("0000010000011111","1100000000100010"),
								 ("0000010000000110","1100000000100000"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001111010100","1100000000011101"),
								 ("0000001110111011","1100000000011100"),
								 ("0000001110100001","1100000000011010"),
								 ("0000001110001000","1100000000011001"),
								 ("0000001101101111","1100000000011000"),
								 ("0000001101010110","1100000000010110"),
								 ("0000001100111101","1100000000010101"),
								 ("0000001100100100","1100000000010100"),
								 ("0000001100001011","1100000000010011"),
								 ("0000001011110010","1100000000010001"),
								 ("0000001011011001","1100000000010000"),
								 ("0000001011000000","1100000000001111"),
								 ("0000001010100110","1100000000001110"),
								 ("0000001010001101","1100000000001101"),
								 ("0000001001110100","1100000000001100"),
								 ("0000001001011011","1100000000001011"),
								 ("0000001001000010","1100000000001010"),
								 ("0000001000101001","1100000000001001"),
								 ("0000001000010000","1100000000001001"),
								 ("0000000111110111","1100000000001000"),
								 ("0000000111011101","1100000000000111"),
								 ("0000000111000100","1100000000000110"),
								 ("0000000110101011","1100000000000110"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000101111001","1100000000000100"),
								 ("0000000101100000","1100000000000100"),
								 ("0000000101000111","1100000000000011"),
								 ("0000000100101110","1100000000000011"),
								 ("0000000100010100","1100000000000010"),
								 ("0000000011111011","1100000000000010"),
								 ("0000000011100010","1100000000000010"),
								 ("0000000011001001","1100000000000001"),
								 ("0000000010110000","1100000000000001"),
								 ("0000000010010111","1100000000000001"),
								 ("0000000001111110","1100000000000000"),
								 ("0000000001100101","1100000000000000"),
								 ("0000000001001011","1100000000000000"),
								 ("0000000000110010","1100000000000000"),
								 ("0000000000011001","1100000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","1111111110110101"),
								 ("0011111111111111","1111111101101001"),
								 ("0011111111111110","1111111100011110"),
								 ("0011111111111101","1111111011010010"),
								 ("0011111111111100","1111111010000111"),
								 ("0011111111111010","1111111000111100"),
								 ("0011111111110111","1111110111110000"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111110010","1111110101011010"),
								 ("0011111111101111","1111110100001110"),
								 ("0011111111101011","1111110011000011"),
								 ("0011111111100111","1111110001111000"),
								 ("0011111111100011","1111110000101100"),
								 ("0011111111011110","1111101111100001"),
								 ("0011111111011001","1111101110010110"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111111001110","1111101100000000"),
								 ("0011111111001000","1111101010110100"),
								 ("0011111111000001","1111101001101001"),
								 ("0011111110111011","1111101000011110"),
								 ("0011111110110100","1111100111010011"),
								 ("0011111110101100","1111100110001000"),
								 ("0011111110100100","1111100100111101"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111110010100","1111100010100111"),
								 ("0011111110001011","1111100001011100"),
								 ("0011111110000010","1111100000010001"),
								 ("0011111101111000","1111011111000111"),
								 ("0011111101101110","1111011101111100"),
								 ("0011111101100100","1111011100110001"),
								 ("0011111101011010","1111011011100111"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111101000011","1111011001010001"),
								 ("0011111100111000","1111011000000111"),
								 ("0011111100101100","1111010110111100"),
								 ("0011111100100000","1111010101110010"),
								 ("0011111100010011","1111010100101000"),
								 ("0011111100000110","1111010011011101"),
								 ("0011111011111001","1111010010010011"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111011011101","1111001111111111"),
								 ("0011111011001111","1111001110110101"),
								 ("0011111011000000","1111001101101011"),
								 ("0011111010110001","1111001100100001"),
								 ("0011111010100010","1111001011010111"),
								 ("0011111010010010","1111001010001110"),
								 ("0011111010000010","1111001001000100"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111001100001","1111000110110001"),
								 ("0011111001010000","1111000101100111"),
								 ("0011111000111111","1111000100011110"),
								 ("0011111000101101","1111000011010101"),
								 ("0011111000011011","1111000010001011"),
								 ("0011111000001001","1111000001000010"),
								 ("0011110111110110","1110111111111001"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110111010000","1110111101100111"),
								 ("0011110110111100","1110111100011111"),
								 ("0011110110101000","1110111011010110"),
								 ("0011110110010011","1110111010001101"),
								 ("0011110101111111","1110111001000101"),
								 ("0011110101101010","1110110111111100"),
								 ("0011110101010100","1110110110110100"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110100101000","1110110100100100"),
								 ("0011110100010010","1110110011011100"),
								 ("0011110011111011","1110110010010100"),
								 ("0011110011100100","1110110001001100"),
								 ("0011110011001101","1110110000000101"),
								 ("0011110010110101","1110101110111101"),
								 ("0011110010011101","1110101101110101"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110001101100","1110101011100111"),
								 ("0011110001010011","1110101010100000"),
								 ("0011110000111010","1110101001011001"),
								 ("0011110000100000","1110101000010010"),
								 ("0011110000000110","1110100111001011"),
								 ("0011101111101100","1110100110000100"),
								 ("0011101111010001","1110100100111110"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101110011011","1110100010110001"),
								 ("0011101101111111","1110100001101011"),
								 ("0011101101100011","1110100000100101"),
								 ("0011101101000111","1110011111011111"),
								 ("0011101100101010","1110011110011001"),
								 ("0011101100001110","1110011101010100"),
								 ("0011101011110000","1110011100001110"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101010110101","1110011010000100"),
								 ("0011101010010111","1110011000111111"),
								 ("0011101001111000","1110010111111010"),
								 ("0011101001011001","1110010110110101"),
								 ("0011101000111010","1110010101110000"),
								 ("0011101000011011","1110010100101100"),
								 ("0011100111111011","1110010011100111"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100110111011","1110010001011111"),
								 ("0011100110011010","1110010000011011"),
								 ("0011100101111001","1110001111010111"),
								 ("0011100101011000","1110001110010100"),
								 ("0011100100110110","1110001101010000"),
								 ("0011100100010100","1110001100001101"),
								 ("0011100011110010","1110001011001010"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100010101100","1110001001000100"),
								 ("0011100010001001","1110001000000001"),
								 ("0011100001100110","1110000110111110"),
								 ("0011100001000010","1110000101111100"),
								 ("0011100000011110","1110000100111010"),
								 ("0011011111111001","1110000011111000"),
								 ("0011011111010101","1110000010110110"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011110001010","1110000000110011"),
								 ("0011011101100101","1101111111110001"),
								 ("0011011100111111","1101111110110000"),
								 ("0011011100011000","1101111101101111"),
								 ("0011011011110010","1101111100101111"),
								 ("0011011011001011","1101111011101110"),
								 ("0011011010100100","1101111010101101"),
								 ("0011011001111101","1101111001101101"),
								 ("0011011001010101","1101111000101101"),
								 ("0011011000101101","1101110111101101"),
								 ("0011011000000101","1101110110101101"),
								 ("0011010111011100","1101110101101110"),
								 ("0011010110110011","1101110100101110"),
								 ("0011010110001010","1101110011101111"),
								 ("0011010101100001","1101110010110000"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010100001101","1101110000110011"),
								 ("0011010011100010","1101101111110101"),
								 ("0011010010111000","1101101110110110"),
								 ("0011010010001101","1101101101111000"),
								 ("0011010001100010","1101101100111011"),
								 ("0011010000110110","1101101011111101"),
								 ("0011010000001011","1101101010111111"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001110110010","1101101001000101"),
								 ("0011001110000110","1101101000001000"),
								 ("0011001101011001","1101100111001100"),
								 ("0011001100101100","1101100110001111"),
								 ("0011001011111110","1101100101010011"),
								 ("0011001011010000","1101100100010111"),
								 ("0011001010100011","1101100011011100"),
								 ("0011001001110100","1101100010100000"),
								 ("0011001001000110","1101100001100101"),
								 ("0011001000010111","1101100000101010"),
								 ("0011000111101000","1101011111101111"),
								 ("0011000110111001","1101011110110100"),
								 ("0011000110001001","1101011101111010"),
								 ("0011000101011001","1101011100111111"),
								 ("0011000100101001","1101011100000101"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000011001000","1101011010010010"),
								 ("0011000010010111","1101011001011001"),
								 ("0011000001100110","1101011000011111"),
								 ("0011000000110100","1101010111100110"),
								 ("0011000000000010","1101010110101110"),
								 ("0010111111010000","1101010101110101"),
								 ("0010111110011110","1101010100111101"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111100111001","1101010011001101"),
								 ("0010111100000110","1101010010010110"),
								 ("0010111011010011","1101010001011111"),
								 ("0010111010011111","1101010000101000"),
								 ("0010111001101011","1101001111110001"),
								 ("0010111000110111","1101001110111010"),
								 ("0010111000000011","1101001110000100"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110110011010","1101001100011000"),
								 ("0010110101100101","1101001011100010"),
								 ("0010110100101111","1101001010101101"),
								 ("0010110011111010","1101001001111000"),
								 ("0010110011000100","1101001001000011"),
								 ("0010110010001110","1101001000001110"),
								 ("0010110001011000","1101000111011010"),
								 ("0010110000100001","1101000110100110"),
								 ("0010101111101011","1101000101110010"),
								 ("0010101110110100","1101000100111110"),
								 ("0010101101111101","1101000100001011"),
								 ("0010101101000101","1101000011011000"),
								 ("0010101100001101","1101000010100101"),
								 ("0010101011010110","1101000001110011"),
								 ("0010101010011101","1101000001000000"),
								 ("0010101001100101","1101000000001110"),
								 ("0010101000101100","1100111111011100"),
								 ("0010100111110100","1100111110101011"),
								 ("0010100110111011","1100111101111001"),
								 ("0010100110000001","1100111101001000"),
								 ("0010100101001000","1100111100011000"),
								 ("0010100100001110","1100111011100111"),
								 ("0010100011010100","1100111010110111"),
								 ("0010100010011010","1100111010000111"),
								 ("0010100001100000","1100111001010111"),
								 ("0010100000100101","1100111000101000"),
								 ("0010011111101010","1100110111111001"),
								 ("0010011110101111","1100110111001010"),
								 ("0010011101110100","1100110110011011"),
								 ("0010011100111000","1100110101101101"),
								 ("0010011011111101","1100110100111111"),
								 ("0010011011000001","1100110100010001"),
								 ("0010011010000101","1100110011100011"),
								 ("0010011001001000","1100110010110110"),
								 ("0010011000001100","1100110010001001"),
								 ("0010010111001111","1100110001011101"),
								 ("0010010110010010","1100110000110000"),
								 ("0010010101010101","1100110000000100"),
								 ("0010010100011000","1100101111011000"),
								 ("0010010011011010","1100101110101101"),
								 ("0010010010011100","1100101110000001"),
								 ("0010010001011110","1100101101010110"),
								 ("0010010000100000","1100101100101100"),
								 ("0010001111100010","1100101100000001"),
								 ("0010001110100011","1100101011010111"),
								 ("0010001101100101","1100101010101101"),
								 ("0010001100100110","1100101010000100"),
								 ("0010001011100111","1100101001011011"),
								 ("0010001010100111","1100101000110010"),
								 ("0010001001101000","1100101000001001"),
								 ("0010001000101000","1100100111100000"),
								 ("0010000111101000","1100100110111000"),
								 ("0010000110101000","1100100110010001"),
								 ("0010000101101000","1100100101101001"),
								 ("0010000100101000","1100100101000010"),
								 ("0010000011100111","1100100100011011"),
								 ("0010000010100110","1100100011110100"),
								 ("0010000001100101","1100100011001110"),
								 ("0010000000100100","1100100010101000"),
								 ("0001111111100011","1100100010000010"),
								 ("0001111110100010","1100100001011101"),
								 ("0001111101100000","1100100000111000"),
								 ("0001111100011110","1100100000010011"),
								 ("0001111011011100","1100011111101110"),
								 ("0001111010011010","1100011111001010"),
								 ("0001111001011000","1100011110100110"),
								 ("0001111000010101","1100011110000011"),
								 ("0001110111010011","1100011101011111"),
								 ("0001110110010000","1100011100111101"),
								 ("0001110101001101","1100011100011010"),
								 ("0001110100001010","1100011011110111"),
								 ("0001110011000110","1100011011010101"),
								 ("0001110010000011","1100011010110100"),
								 ("0001110000111111","1100011010010010"),
								 ("0001101111111100","1100011001110001"),
								 ("0001101110111000","1100011001010000"),
								 ("0001101101110100","1100011000110000"),
								 ("0001101100110000","1100011000010000"),
								 ("0001101011101011","1100010111110000"),
								 ("0001101010100111","1100010111010000"),
								 ("0001101001100010","1100010110110001"),
								 ("0001101000011101","1100010110010010"),
								 ("0001100111011000","1100010101110011"),
								 ("0001100110010011","1100010101010101"),
								 ("0001100101001110","1100010100110111"),
								 ("0001100100001001","1100010100011010"),
								 ("0001100011000011","1100010011111100"),
								 ("0001100001111110","1100010011011111"),
								 ("0001100000111000","1100010011000010"),
								 ("0001011111110010","1100010010100110"),
								 ("0001011110101100","1100010010001010"),
								 ("0001011101100110","1100010001101110"),
								 ("0001011100100000","1100010001010011"),
								 ("0001011011011010","1100010000111000"),
								 ("0001011010010011","1100010000011101"),
								 ("0001011001001100","1100010000000011"),
								 ("0001011000000110","1100001111101001"),
								 ("0001010110111111","1100001111001111"),
								 ("0001010101111000","1100001110110101"),
								 ("0001010100110001","1100001110011100"),
								 ("0001010011101010","1100001110000011"),
								 ("0001010010100010","1100001101101011"),
								 ("0001010001011011","1100001101010011"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001111001100","1100001100100011"),
								 ("0001001110000100","1100001100001100"),
								 ("0001001100111100","1100001011110101"),
								 ("0001001011110100","1100001011011111"),
								 ("0001001010101100","1100001011001001"),
								 ("0001001001100100","1100001010110011"),
								 ("0001001000011100","1100001010011101"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000110001011","1100001001110011"),
								 ("0001000101000010","1100001001011111"),
								 ("0001000011111010","1100001001001011"),
								 ("0001000010110001","1100001000110111"),
								 ("0001000001101000","1100001000100011"),
								 ("0001000000011111","1100001000010000"),
								 ("0000111111010110","1100000111111101"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111101000100","1100000111011001"),
								 ("0000111011111011","1100000111000111"),
								 ("0000111010110001","1100000110110110"),
								 ("0000111001101000","1100000110100100"),
								 ("0000111000011110","1100000110010100"),
								 ("0000110111010101","1100000110000011"),
								 ("0000110110001011","1100000101110011"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110011111000","1100000101010100"),
								 ("0000110010101110","1100000101000101"),
								 ("0000110001100100","1100000100110110"),
								 ("0000110000011010","1100000100101000"),
								 ("0000101111010000","1100000100011001"),
								 ("0000101110000101","1100000100001100"),
								 ("0000101100111011","1100000011111110"),
								 ("0000101011110001","1100000011110001"),
								 ("0000101010100111","1100000011100100"),
								 ("0000101001011100","1100000011011000"),
								 ("0000101000010010","1100000011001100"),
								 ("0000100111000111","1100000011000000"),
								 ("0000100101111101","1100000010110101"),
								 ("0000100100110010","1100000010101010"),
								 ("0000100011101000","1100000010011111"),
								 ("0000100010011101","1100000010010101"),
								 ("0000100001010010","1100000010001011"),
								 ("0000100000000111","1100000010000001"),
								 ("0000011110111101","1100000001111000"),
								 ("0000011101110010","1100000001101111"),
								 ("0000011100100111","1100000001100111"),
								 ("0000011011011100","1100000001011110"),
								 ("0000011010010001","1100000001010110"),
								 ("0000011001000110","1100000001001111"),
								 ("0000010111111011","1100000001001000"),
								 ("0000010110110000","1100000001000001"),
								 ("0000010101100101","1100000000111010"),
								 ("0000010100011010","1100000000110100"),
								 ("0000010011001110","1100000000101110"),
								 ("0000010010000011","1100000000101001"),
								 ("0000010000111000","1100000000100100"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001110100001","1100000000011010"),
								 ("0000001101010110","1100000000010110"),
								 ("0000001100001011","1100000000010011"),
								 ("0000001011000000","1100000000001111"),
								 ("0000001001110100","1100000000001100"),
								 ("0000001000101001","1100000000001001"),
								 ("0000000111011101","1100000000000111"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000101000111","1100000000000011"),
								 ("0000000011111011","1100000000000010"),
								 ("0000000010110000","1100000000000001"),
								 ("0000000001100101","1100000000000000"),
								 ("0000000000011001","1100000000000000"),
								 ("1111111111001110","1100000000000000"),
								 ("1111111110000010","1100000000000000"),
								 ("1111111100110111","1100000000000001"),
								 ("1111111011101100","1100000000000010"),
								 ("1111111010100000","1100000000000100"),
								 ("1111111001010101","1100000000000110"),
								 ("1111111000001001","1100000000001000"),
								 ("1111110110111110","1100000000001010"),
								 ("1111110101110011","1100000000001101"),
								 ("1111110100100111","1100000000010000"),
								 ("1111110011011100","1100000000010100"),
								 ("1111110010010001","1100000000011000"),
								 ("1111110001000101","1100000000011100"),
								 ("1111101111111010","1100000000100000"),
								 ("1111101110101111","1100000000100101"),
								 ("1111101101100100","1100000000101011"),
								 ("1111101100011001","1100000000110000"),
								 ("1111101011001101","1100000000110110"),
								 ("1111101010000010","1100000000111100"),
								 ("1111101000110111","1100000001000011"),
								 ("1111100111101100","1100000001001010"),
								 ("1111100110100001","1100000001010001"),
								 ("1111100101010110","1100000001011001"),
								 ("1111100100001011","1100000001100001"),
								 ("1111100011000000","1100000001101001"),
								 ("1111100001110101","1100000001110010"),
								 ("1111100000101010","1100000001111011"),
								 ("1111011111100000","1100000010000101"),
								 ("1111011110010101","1100000010001110"),
								 ("1111011101001010","1100000010011000"),
								 ("1111011011111111","1100000010100011"),
								 ("1111011010110101","1100000010101110"),
								 ("1111011001101010","1100000010111001"),
								 ("1111011000100000","1100000011000100"),
								 ("1111010111010101","1100000011010000"),
								 ("1111010110001011","1100000011011100"),
								 ("1111010101000000","1100000011101001"),
								 ("1111010011110110","1100000011110110"),
								 ("1111010010101100","1100000100000011"),
								 ("1111010001100010","1100000100010000"),
								 ("1111010000011000","1100000100011110"),
								 ("1111001111001110","1100000100101100"),
								 ("1111001110000100","1100000100111011"),
								 ("1111001100111010","1100000101001010"),
								 ("1111001011110000","1100000101011001"),
								 ("1111001010100110","1100000101101000"),
								 ("1111001001011100","1100000101111000"),
								 ("1111001000010011","1100000110001001"),
								 ("1111000111001001","1100000110011001"),
								 ("1111000110000000","1100000110101010"),
								 ("1111000100110110","1100000110111011"),
								 ("1111000011101101","1100000111001101"),
								 ("1111000010100100","1100000111011111"),
								 ("1111000001011011","1100000111110001"),
								 ("1111000000010010","1100001000000100"),
								 ("1110111111001001","1100001000010111"),
								 ("1110111110000000","1100001000101010"),
								 ("1110111100110111","1100001000111110"),
								 ("1110111011101110","1100001001010001"),
								 ("1110111010100110","1100001001100110"),
								 ("1110111001011101","1100001001111010"),
								 ("1110111000010101","1100001010001111"),
								 ("1110110111001100","1100001010100101"),
								 ("1110110110000100","1100001010111010"),
								 ("1110110100111100","1100001011010000"),
								 ("1110110011110100","1100001011100110"),
								 ("1110110010101100","1100001011111101"),
								 ("1110110001100100","1100001100010100"),
								 ("1110110000011100","1100001100101011"),
								 ("1110101111010101","1100001101000011"),
								 ("1110101110001101","1100001101011011"),
								 ("1110101101000110","1100001101110011"),
								 ("1110101011111111","1100001110001100"),
								 ("1110101010110111","1100001110100101"),
								 ("1110101001110000","1100001110111110"),
								 ("1110101000101001","1100001111010111"),
								 ("1110100111100011","1100001111110001"),
								 ("1110100110011100","1100010000001011"),
								 ("1110100101010101","1100010000100110"),
								 ("1110100100001111","1100010001000001"),
								 ("1110100011001001","1100010001011100"),
								 ("1110100010000010","1100010001111000"),
								 ("1110100000111100","1100010010010011"),
								 ("1110011111110110","1100010010110000"),
								 ("1110011110110001","1100010011001100"),
								 ("1110011101101011","1100010011101001"),
								 ("1110011100100101","1100010100000110"),
								 ("1110011011100000","1100010100100011"),
								 ("1110011010011011","1100010101000001"),
								 ("1110011001010110","1100010101011111"),
								 ("1110011000010001","1100010101111110"),
								 ("1110010111001100","1100010110011100"),
								 ("1110010110000111","1100010110111011"),
								 ("1110010101000010","1100010111011011"),
								 ("1110010011111110","1100010111111010"),
								 ("1110010010111010","1100011000011010"),
								 ("1110010001110110","1100011000111011"),
								 ("1110010000110010","1100011001011011"),
								 ("1110001111101110","1100011001111100"),
								 ("1110001110101010","1100011010011101"),
								 ("1110001101100111","1100011010111111"),
								 ("1110001100100011","1100011011100001"),
								 ("1110001011100000","1100011100000011"),
								 ("1110001010011101","1100011100100101"),
								 ("1110001001011010","1100011101001000"),
								 ("1110001000010111","1100011101101011"),
								 ("1110000111010101","1100011110001111"),
								 ("1110000110010010","1100011110110010"),
								 ("1110000101010000","1100011111010110"),
								 ("1110000100001110","1100011111111011"),
								 ("1110000011001100","1100100000011111"),
								 ("1110000010001010","1100100001000100"),
								 ("1110000001001001","1100100001101001"),
								 ("1110000000000111","1100100010001111"),
								 ("1101111111000110","1100100010110101"),
								 ("1101111110000101","1100100011011011"),
								 ("1101111101000100","1100100100000001"),
								 ("1101111100000011","1100100100101000"),
								 ("1101111011000011","1100100101001111"),
								 ("1101111010000011","1100100101110110"),
								 ("1101111001000010","1100100110011110"),
								 ("1101111000000010","1100100111000110"),
								 ("1101110111000011","1100100111101110"),
								 ("1101110110000011","1100101000010110"),
								 ("1101110101000100","1100101000111111"),
								 ("1101110100000100","1100101001101000"),
								 ("1101110011000101","1100101010010010"),
								 ("1101110010000110","1100101010111011"),
								 ("1101110001001000","1100101011100101"),
								 ("1101110000001001","1100101100001111"),
								 ("1101101111001011","1100101100111010"),
								 ("1101101110001101","1100101101100101"),
								 ("1101101101001111","1100101110010000"),
								 ("1101101100010001","1100101110111011"),
								 ("1101101011010100","1100101111100111"),
								 ("1101101010010111","1100110000010011"),
								 ("1101101001011010","1100110000111111"),
								 ("1101101000011101","1100110001101011"),
								 ("1101100111100000","1100110010011000"),
								 ("1101100110100100","1100110011000101"),
								 ("1101100101100111","1100110011110011"),
								 ("1101100100101011","1100110100100000"),
								 ("1101100011101111","1100110101001110"),
								 ("1101100010110100","1100110101111100"),
								 ("1101100001111000","1100110110101011"),
								 ("1101100000111101","1100110111011001"),
								 ("1101100000000010","1100111000001000"),
								 ("1101011111001000","1100111000111000"),
								 ("1101011110001101","1100111001100111"),
								 ("1101011101010011","1100111010010111"),
								 ("1101011100011001","1100111011000111"),
								 ("1101011011011111","1100111011110111"),
								 ("1101011010100101","1100111100101000"),
								 ("1101011001101100","1100111101011001"),
								 ("1101011000110010","1100111110001010"),
								 ("1101010111111001","1100111110111011"),
								 ("1101010111000001","1100111111101101"),
								 ("1101010110001000","1101000000011111"),
								 ("1101010101010000","1101000001010001"),
								 ("1101010100011000","1101000010000011"),
								 ("1101010011100000","1101000010110110"),
								 ("1101010010101000","1101000011101001"),
								 ("1101010001110001","1101000100011100"),
								 ("1101010000111010","1101000101010000"),
								 ("1101010000000011","1101000110000011"),
								 ("1101001111001100","1101000110110111"),
								 ("1101001110010110","1101000111101011"),
								 ("1101001101100000","1101001000100000"),
								 ("1101001100101010","1101001001010101"),
								 ("1101001011110100","1101001010001010"),
								 ("1101001010111111","1101001010111111"),
								 ("1101001010001010","1101001011110100"),
								 ("1101001001010101","1101001100101010"),
								 ("1101001000100000","1101001101100000"),
								 ("1101000111101011","1101001110010110"),
								 ("1101000110110111","1101001111001100"),
								 ("1101000110000011","1101010000000011"),
								 ("1101000101010000","1101010000111010"),
								 ("1101000100011100","1101010001110001"),
								 ("1101000011101001","1101010010101000"),
								 ("1101000010110110","1101010011100000"),
								 ("1101000010000011","1101010100011000"),
								 ("1101000001010001","1101010101010000"),
								 ("1101000000011111","1101010110001000"),
								 ("1100111111101101","1101010111000001"),
								 ("1100111110111011","1101010111111001"),
								 ("1100111110001010","1101011000110010"),
								 ("1100111101011001","1101011001101100"),
								 ("1100111100101000","1101011010100101"),
								 ("1100111011110111","1101011011011111"),
								 ("1100111011000111","1101011100011001"),
								 ("1100111010010111","1101011101010011"),
								 ("1100111001100111","1101011110001101"),
								 ("1100111000111000","1101011111001000"),
								 ("1100111000001000","1101100000000010"),
								 ("1100110111011001","1101100000111101"),
								 ("1100110110101011","1101100001111000"),
								 ("1100110101111100","1101100010110100"),
								 ("1100110101001110","1101100011101111"),
								 ("1100110100100000","1101100100101011"),
								 ("1100110011110011","1101100101100111"),
								 ("1100110011000101","1101100110100100"),
								 ("1100110010011000","1101100111100000"),
								 ("1100110001101011","1101101000011101"),
								 ("1100110000111111","1101101001011010"),
								 ("1100110000010011","1101101010010111"),
								 ("1100101111100111","1101101011010100"),
								 ("1100101110111011","1101101100010001"),
								 ("1100101110010000","1101101101001111"),
								 ("1100101101100101","1101101110001101"),
								 ("1100101100111010","1101101111001011"),
								 ("1100101100001111","1101110000001001"),
								 ("1100101011100101","1101110001001000"),
								 ("1100101010111011","1101110010000110"),
								 ("1100101010010010","1101110011000101"),
								 ("1100101001101000","1101110100000100"),
								 ("1100101000111111","1101110101000100"),
								 ("1100101000010110","1101110110000011"),
								 ("1100100111101110","1101110111000011"),
								 ("1100100111000110","1101111000000010"),
								 ("1100100110011110","1101111001000010"),
								 ("1100100101110110","1101111010000011"),
								 ("1100100101001111","1101111011000011"),
								 ("1100100100101000","1101111100000011"),
								 ("1100100100000001","1101111101000100"),
								 ("1100100011011011","1101111110000101"),
								 ("1100100010110101","1101111111000110"),
								 ("1100100010001111","1110000000000111"),
								 ("1100100001101001","1110000001001001"),
								 ("1100100001000100","1110000010001010"),
								 ("1100100000011111","1110000011001100"),
								 ("1100011111111011","1110000100001110"),
								 ("1100011111010110","1110000101010000"),
								 ("1100011110110010","1110000110010010"),
								 ("1100011110001111","1110000111010101"),
								 ("1100011101101011","1110001000010111"),
								 ("1100011101001000","1110001001011010"),
								 ("1100011100100101","1110001010011101"),
								 ("1100011100000011","1110001011100000"),
								 ("1100011011100001","1110001100100011"),
								 ("1100011010111111","1110001101100111"),
								 ("1100011010011101","1110001110101010"),
								 ("1100011001111100","1110001111101110"),
								 ("1100011001011011","1110010000110010"),
								 ("1100011000111011","1110010001110110"),
								 ("1100011000011010","1110010010111010"),
								 ("1100010111111010","1110010011111110"),
								 ("1100010111011011","1110010101000010"),
								 ("1100010110111011","1110010110000111"),
								 ("1100010110011100","1110010111001100"),
								 ("1100010101111110","1110011000010001"),
								 ("1100010101011111","1110011001010110"),
								 ("1100010101000001","1110011010011011"),
								 ("1100010100100011","1110011011100000"),
								 ("1100010100000110","1110011100100101"),
								 ("1100010011101001","1110011101101011"),
								 ("1100010011001100","1110011110110001"),
								 ("1100010010110000","1110011111110110"),
								 ("1100010010010011","1110100000111100"),
								 ("1100010001111000","1110100010000010"),
								 ("1100010001011100","1110100011001001"),
								 ("1100010001000001","1110100100001111"),
								 ("1100010000100110","1110100101010101"),
								 ("1100010000001011","1110100110011100"),
								 ("1100001111110001","1110100111100011"),
								 ("1100001111010111","1110101000101001"),
								 ("1100001110111110","1110101001110000"),
								 ("1100001110100101","1110101010110111"),
								 ("1100001110001100","1110101011111111"),
								 ("1100001101110011","1110101101000110"),
								 ("1100001101011011","1110101110001101"),
								 ("1100001101000011","1110101111010101"),
								 ("1100001100101011","1110110000011100"),
								 ("1100001100010100","1110110001100100"),
								 ("1100001011111101","1110110010101100"),
								 ("1100001011100110","1110110011110100"),
								 ("1100001011010000","1110110100111100"),
								 ("1100001010111010","1110110110000100"),
								 ("1100001010100101","1110110111001100"),
								 ("1100001010001111","1110111000010101"),
								 ("1100001001111010","1110111001011101"),
								 ("1100001001100110","1110111010100110"),
								 ("1100001001010001","1110111011101110"),
								 ("1100001000111110","1110111100110111"),
								 ("1100001000101010","1110111110000000"),
								 ("1100001000010111","1110111111001001"),
								 ("1100001000000100","1111000000010010"),
								 ("1100000111110001","1111000001011011"),
								 ("1100000111011111","1111000010100100"),
								 ("1100000111001101","1111000011101101"),
								 ("1100000110111011","1111000100110110"),
								 ("1100000110101010","1111000110000000"),
								 ("1100000110011001","1111000111001001"),
								 ("1100000110001001","1111001000010011"),
								 ("1100000101111000","1111001001011100"),
								 ("1100000101101000","1111001010100110"),
								 ("1100000101011001","1111001011110000"),
								 ("1100000101001010","1111001100111010"),
								 ("1100000100111011","1111001110000100"),
								 ("1100000100101100","1111001111001110"),
								 ("1100000100011110","1111010000011000"),
								 ("1100000100010000","1111010001100010"),
								 ("1100000100000011","1111010010101100"),
								 ("1100000011110110","1111010011110110"),
								 ("1100000011101001","1111010101000000"),
								 ("1100000011011100","1111010110001011"),
								 ("1100000011010000","1111010111010101"),
								 ("1100000011000100","1111011000100000"),
								 ("1100000010111001","1111011001101010"),
								 ("1100000010101110","1111011010110101"),
								 ("1100000010100011","1111011011111111"),
								 ("1100000010011000","1111011101001010"),
								 ("1100000010001110","1111011110010101"),
								 ("1100000010000101","1111011111100000"),
								 ("1100000001111011","1111100000101010"),
								 ("1100000001110010","1111100001110101"),
								 ("1100000001101001","1111100011000000"),
								 ("1100000001100001","1111100100001011"),
								 ("1100000001011001","1111100101010110"),
								 ("1100000001010001","1111100110100001"),
								 ("1100000001001010","1111100111101100"),
								 ("1100000001000011","1111101000110111"),
								 ("1100000000111100","1111101010000010"),
								 ("1100000000110110","1111101011001101"),
								 ("1100000000110000","1111101100011001"),
								 ("1100000000101011","1111101101100100"),
								 ("1100000000100101","1111101110101111"),
								 ("1100000000100000","1111101111111010"),
								 ("1100000000011100","1111110001000101"),
								 ("1100000000011000","1111110010010001"),
								 ("1100000000010100","1111110011011100"),
								 ("1100000000010000","1111110100100111"),
								 ("1100000000001101","1111110101110011"),
								 ("1100000000001010","1111110110111110"),
								 ("1100000000001000","1111111000001001"),
								 ("1100000000000110","1111111001010101"),
								 ("1100000000000100","1111111010100000"),
								 ("1100000000000010","1111111011101100"),
								 ("1100000000000001","1111111100110111"),
								 ("1100000000000000","1111111110000010"),
								 ("1100000000000000","1111111111001110"),
								 ("1100000000000000","0000000000011001"),
								 ("1100000000000000","0000000001100101"),
								 ("1100000000000001","0000000010110000"),
								 ("1100000000000010","0000000011111011"),
								 ("1100000000000011","0000000101000111"),
								 ("1100000000000101","0000000110010010"),
								 ("1100000000000111","0000000111011101"),
								 ("1100000000001001","0000001000101001"),
								 ("1100000000001100","0000001001110100"),
								 ("1100000000001111","0000001011000000"),
								 ("1100000000010011","0000001100001011"),
								 ("1100000000010110","0000001101010110"),
								 ("1100000000011010","0000001110100001"),
								 ("1100000000011111","0000001111101101"),
								 ("1100000000100100","0000010000111000"),
								 ("1100000000101001","0000010010000011"),
								 ("1100000000101110","0000010011001110"),
								 ("1100000000110100","0000010100011010"),
								 ("1100000000111010","0000010101100101"),
								 ("1100000001000001","0000010110110000"),
								 ("1100000001001000","0000010111111011"),
								 ("1100000001001111","0000011001000110"),
								 ("1100000001010110","0000011010010001"),
								 ("1100000001011110","0000011011011100"),
								 ("1100000001100111","0000011100100111"),
								 ("1100000001101111","0000011101110010"),
								 ("1100000001111000","0000011110111101"),
								 ("1100000010000001","0000100000000111"),
								 ("1100000010001011","0000100001010010"),
								 ("1100000010010101","0000100010011101"),
								 ("1100000010011111","0000100011101000"),
								 ("1100000010101010","0000100100110010"),
								 ("1100000010110101","0000100101111101"),
								 ("1100000011000000","0000100111000111"),
								 ("1100000011001100","0000101000010010"),
								 ("1100000011011000","0000101001011100"),
								 ("1100000011100100","0000101010100111"),
								 ("1100000011110001","0000101011110001"),
								 ("1100000011111110","0000101100111011"),
								 ("1100000100001100","0000101110000101"),
								 ("1100000100011001","0000101111010000"),
								 ("1100000100101000","0000110000011010"),
								 ("1100000100110110","0000110001100100"),
								 ("1100000101000101","0000110010101110"),
								 ("1100000101010100","0000110011111000"),
								 ("1100000101100011","0000110101000001"),
								 ("1100000101110011","0000110110001011"),
								 ("1100000110000011","0000110111010101"),
								 ("1100000110010100","0000111000011110"),
								 ("1100000110100100","0000111001101000"),
								 ("1100000110110110","0000111010110001"),
								 ("1100000111000111","0000111011111011"),
								 ("1100000111011001","0000111101000100"),
								 ("1100000111101011","0000111110001101"),
								 ("1100000111111101","0000111111010110"),
								 ("1100001000010000","0001000000011111"),
								 ("1100001000100011","0001000001101000"),
								 ("1100001000110111","0001000010110001"),
								 ("1100001001001011","0001000011111010"),
								 ("1100001001011111","0001000101000010"),
								 ("1100001001110011","0001000110001011"),
								 ("1100001010001000","0001000111010011"),
								 ("1100001010011101","0001001000011100"),
								 ("1100001010110011","0001001001100100"),
								 ("1100001011001001","0001001010101100"),
								 ("1100001011011111","0001001011110100"),
								 ("1100001011110101","0001001100111100"),
								 ("1100001100001100","0001001110000100"),
								 ("1100001100100011","0001001111001100"),
								 ("1100001100111011","0001010000010011"),
								 ("1100001101010011","0001010001011011"),
								 ("1100001101101011","0001010010100010"),
								 ("1100001110000011","0001010011101010"),
								 ("1100001110011100","0001010100110001"),
								 ("1100001110110101","0001010101111000"),
								 ("1100001111001111","0001010110111111"),
								 ("1100001111101001","0001011000000110"),
								 ("1100010000000011","0001011001001100"),
								 ("1100010000011101","0001011010010011"),
								 ("1100010000111000","0001011011011010"),
								 ("1100010001010011","0001011100100000"),
								 ("1100010001101110","0001011101100110"),
								 ("1100010010001010","0001011110101100"),
								 ("1100010010100110","0001011111110010"),
								 ("1100010011000010","0001100000111000"),
								 ("1100010011011111","0001100001111110"),
								 ("1100010011111100","0001100011000011"),
								 ("1100010100011010","0001100100001001"),
								 ("1100010100110111","0001100101001110"),
								 ("1100010101010101","0001100110010011"),
								 ("1100010101110011","0001100111011000"),
								 ("1100010110010010","0001101000011101"),
								 ("1100010110110001","0001101001100010"),
								 ("1100010111010000","0001101010100111"),
								 ("1100010111110000","0001101011101011"),
								 ("1100011000010000","0001101100110000"),
								 ("1100011000110000","0001101101110100"),
								 ("1100011001010000","0001101110111000"),
								 ("1100011001110001","0001101111111100"),
								 ("1100011010010010","0001110000111111"),
								 ("1100011010110100","0001110010000011"),
								 ("1100011011010101","0001110011000110"),
								 ("1100011011110111","0001110100001010"),
								 ("1100011100011010","0001110101001101"),
								 ("1100011100111101","0001110110010000"),
								 ("1100011101011111","0001110111010011"),
								 ("1100011110000011","0001111000010101"),
								 ("1100011110100110","0001111001011000"),
								 ("1100011111001010","0001111010011010"),
								 ("1100011111101110","0001111011011100"),
								 ("1100100000010011","0001111100011110"),
								 ("1100100000111000","0001111101100000"),
								 ("1100100001011101","0001111110100010"),
								 ("1100100010000010","0001111111100011"),
								 ("1100100010101000","0010000000100100"),
								 ("1100100011001110","0010000001100101"),
								 ("1100100011110100","0010000010100110"),
								 ("1100100100011011","0010000011100111"),
								 ("1100100101000010","0010000100101000"),
								 ("1100100101101001","0010000101101000"),
								 ("1100100110010001","0010000110101000"),
								 ("1100100110111000","0010000111101000"),
								 ("1100100111100000","0010001000101000"),
								 ("1100101000001001","0010001001101000"),
								 ("1100101000110010","0010001010100111"),
								 ("1100101001011011","0010001011100111"),
								 ("1100101010000100","0010001100100110"),
								 ("1100101010101101","0010001101100101"),
								 ("1100101011010111","0010001110100011"),
								 ("1100101100000001","0010001111100010"),
								 ("1100101100101100","0010010000100000"),
								 ("1100101101010110","0010010001011110"),
								 ("1100101110000001","0010010010011100"),
								 ("1100101110101101","0010010011011010"),
								 ("1100101111011000","0010010100011000"),
								 ("1100110000000100","0010010101010101"),
								 ("1100110000110000","0010010110010010"),
								 ("1100110001011101","0010010111001111"),
								 ("1100110010001001","0010011000001100"),
								 ("1100110010110110","0010011001001000"),
								 ("1100110011100011","0010011010000101"),
								 ("1100110100010001","0010011011000001"),
								 ("1100110100111111","0010011011111101"),
								 ("1100110101101101","0010011100111000"),
								 ("1100110110011011","0010011101110100"),
								 ("1100110111001010","0010011110101111"),
								 ("1100110111111001","0010011111101010"),
								 ("1100111000101000","0010100000100101"),
								 ("1100111001010111","0010100001100000"),
								 ("1100111010000111","0010100010011010"),
								 ("1100111010110111","0010100011010100"),
								 ("1100111011100111","0010100100001110"),
								 ("1100111100011000","0010100101001000"),
								 ("1100111101001000","0010100110000001"),
								 ("1100111101111001","0010100110111011"),
								 ("1100111110101011","0010100111110100"),
								 ("1100111111011100","0010101000101100"),
								 ("1101000000001110","0010101001100101"),
								 ("1101000001000000","0010101010011101"),
								 ("1101000001110011","0010101011010110"),
								 ("1101000010100101","0010101100001101"),
								 ("1101000011011000","0010101101000101"),
								 ("1101000100001011","0010101101111101"),
								 ("1101000100111110","0010101110110100"),
								 ("1101000101110010","0010101111101011"),
								 ("1101000110100110","0010110000100001"),
								 ("1101000111011010","0010110001011000"),
								 ("1101001000001110","0010110010001110"),
								 ("1101001001000011","0010110011000100"),
								 ("1101001001111000","0010110011111010"),
								 ("1101001010101101","0010110100101111"),
								 ("1101001011100010","0010110101100101"),
								 ("1101001100011000","0010110110011010"),
								 ("1101001101001110","0010110111001111"),
								 ("1101001110000100","0010111000000011"),
								 ("1101001110111010","0010111000110111"),
								 ("1101001111110001","0010111001101011"),
								 ("1101010000101000","0010111010011111"),
								 ("1101010001011111","0010111011010011"),
								 ("1101010010010110","0010111100000110"),
								 ("1101010011001101","0010111100111001"),
								 ("1101010100000101","0010111101101100"),
								 ("1101010100111101","0010111110011110"),
								 ("1101010101110101","0010111111010000"),
								 ("1101010110101110","0011000000000010"),
								 ("1101010111100110","0011000000110100"),
								 ("1101011000011111","0011000001100110"),
								 ("1101011001011001","0011000010010111"),
								 ("1101011010010010","0011000011001000"),
								 ("1101011011001011","0011000011111001"),
								 ("1101011100000101","0011000100101001"),
								 ("1101011100111111","0011000101011001"),
								 ("1101011101111010","0011000110001001"),
								 ("1101011110110100","0011000110111001"),
								 ("1101011111101111","0011000111101000"),
								 ("1101100000101010","0011001000010111"),
								 ("1101100001100101","0011001001000110"),
								 ("1101100010100000","0011001001110100"),
								 ("1101100011011100","0011001010100011"),
								 ("1101100100010111","0011001011010000"),
								 ("1101100101010011","0011001011111110"),
								 ("1101100110001111","0011001100101100"),
								 ("1101100111001100","0011001101011001"),
								 ("1101101000001000","0011001110000110"),
								 ("1101101001000101","0011001110110010"),
								 ("1101101010000010","0011001111011111"),
								 ("1101101010111111","0011010000001011"),
								 ("1101101011111101","0011010000110110"),
								 ("1101101100111011","0011010001100010"),
								 ("1101101101111000","0011010010001101"),
								 ("1101101110110110","0011010010111000"),
								 ("1101101111110101","0011010011100010"),
								 ("1101110000110011","0011010100001101"),
								 ("1101110001110010","0011010100110111"),
								 ("1101110010110000","0011010101100001"),
								 ("1101110011101111","0011010110001010"),
								 ("1101110100101110","0011010110110011"),
								 ("1101110101101110","0011010111011100"),
								 ("1101110110101101","0011011000000101"),
								 ("1101110111101101","0011011000101101"),
								 ("1101111000101101","0011011001010101"),
								 ("1101111001101101","0011011001111101"),
								 ("1101111010101101","0011011010100100"),
								 ("1101111011101110","0011011011001011"),
								 ("1101111100101111","0011011011110010"),
								 ("1101111101101111","0011011100011000"),
								 ("1101111110110000","0011011100111111"),
								 ("1101111111110001","0011011101100101"),
								 ("1110000000110011","0011011110001010"),
								 ("1110000001110100","0011011110110000"),
								 ("1110000010110110","0011011111010101"),
								 ("1110000011111000","0011011111111001"),
								 ("1110000100111010","0011100000011110"),
								 ("1110000101111100","0011100001000010"),
								 ("1110000110111110","0011100001100110"),
								 ("1110001000000001","0011100010001001"),
								 ("1110001001000100","0011100010101100"),
								 ("1110001010000111","0011100011001111"),
								 ("1110001011001010","0011100011110010"),
								 ("1110001100001101","0011100100010100"),
								 ("1110001101010000","0011100100110110"),
								 ("1110001110010100","0011100101011000"),
								 ("1110001111010111","0011100101111001"),
								 ("1110010000011011","0011100110011010"),
								 ("1110010001011111","0011100110111011"),
								 ("1110010010100011","0011100111011011"),
								 ("1110010011100111","0011100111111011"),
								 ("1110010100101100","0011101000011011"),
								 ("1110010101110000","0011101000111010"),
								 ("1110010110110101","0011101001011001"),
								 ("1110010111111010","0011101001111000"),
								 ("1110011000111111","0011101010010111"),
								 ("1110011010000100","0011101010110101"),
								 ("1110011011001001","0011101011010011"),
								 ("1110011100001110","0011101011110000"),
								 ("1110011101010100","0011101100001110"),
								 ("1110011110011001","0011101100101010"),
								 ("1110011111011111","0011101101000111"),
								 ("1110100000100101","0011101101100011"),
								 ("1110100001101011","0011101101111111"),
								 ("1110100010110001","0011101110011011"),
								 ("1110100011110111","0011101110110110"),
								 ("1110100100111110","0011101111010001"),
								 ("1110100110000100","0011101111101100"),
								 ("1110100111001011","0011110000000110"),
								 ("1110101000010010","0011110000100000"),
								 ("1110101001011001","0011110000111010"),
								 ("1110101010100000","0011110001010011"),
								 ("1110101011100111","0011110001101100"),
								 ("1110101100101110","0011110010000101"),
								 ("1110101101110101","0011110010011101"),
								 ("1110101110111101","0011110010110101"),
								 ("1110110000000101","0011110011001101"),
								 ("1110110001001100","0011110011100100"),
								 ("1110110010010100","0011110011111011"),
								 ("1110110011011100","0011110100010010"),
								 ("1110110100100100","0011110100101000"),
								 ("1110110101101100","0011110100111111"),
								 ("1110110110110100","0011110101010100"),
								 ("1110110111111100","0011110101101010"),
								 ("1110111001000101","0011110101111111"),
								 ("1110111010001101","0011110110010011"),
								 ("1110111011010110","0011110110101000"),
								 ("1110111100011111","0011110110111100"),
								 ("1110111101100111","0011110111010000"),
								 ("1110111110110000","0011110111100011"),
								 ("1110111111111001","0011110111110110"),
								 ("1111000001000010","0011111000001001"),
								 ("1111000010001011","0011111000011011"),
								 ("1111000011010101","0011111000101101"),
								 ("1111000100011110","0011111000111111"),
								 ("1111000101100111","0011111001010000"),
								 ("1111000110110001","0011111001100001"),
								 ("1111000111111010","0011111001110010"),
								 ("1111001001000100","0011111010000010"),
								 ("1111001010001110","0011111010010010"),
								 ("1111001011010111","0011111010100010"),
								 ("1111001100100001","0011111010110001"),
								 ("1111001101101011","0011111011000000"),
								 ("1111001110110101","0011111011001111"),
								 ("1111001111111111","0011111011011101"),
								 ("1111010001001001","0011111011101011"),
								 ("1111010010010011","0011111011111001"),
								 ("1111010011011101","0011111100000110"),
								 ("1111010100101000","0011111100010011"),
								 ("1111010101110010","0011111100100000"),
								 ("1111010110111100","0011111100101100"),
								 ("1111011000000111","0011111100111000"),
								 ("1111011001010001","0011111101000011"),
								 ("1111011010011100","0011111101001111"),
								 ("1111011011100111","0011111101011010"),
								 ("1111011100110001","0011111101100100"),
								 ("1111011101111100","0011111101101110"),
								 ("1111011111000111","0011111101111000"),
								 ("1111100000010001","0011111110000010"),
								 ("1111100001011100","0011111110001011"),
								 ("1111100010100111","0011111110010100"),
								 ("1111100011110010","0011111110011100"),
								 ("1111100100111101","0011111110100100"),
								 ("1111100110001000","0011111110101100"),
								 ("1111100111010011","0011111110110100"),
								 ("1111101000011110","0011111110111011"),
								 ("1111101001101001","0011111111000001"),
								 ("1111101010110100","0011111111001000"),
								 ("1111101100000000","0011111111001110"),
								 ("1111101101001011","0011111111010100"),
								 ("1111101110010110","0011111111011001"),
								 ("1111101111100001","0011111111011110"),
								 ("1111110000101100","0011111111100011"),
								 ("1111110001111000","0011111111100111"),
								 ("1111110011000011","0011111111101011"),
								 ("1111110100001110","0011111111101111"),
								 ("1111110101011010","0011111111110010"),
								 ("1111110110100101","0011111111110101"),
								 ("1111110111110000","0011111111110111"),
								 ("1111111000111100","0011111111111010"),
								 ("1111111010000111","0011111111111100"),
								 ("1111111011010010","0011111111111101"),
								 ("1111111100011110","0011111111111110"),
								 ("1111111101101001","0011111111111111"),
								 ("1111111110110101","0100000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000")
							   );
begin
	doutr <= std_logic_vector(rom(conv_integer(addr))(0));
	douti <= std_logic_vector(rom(conv_integer(addr))(1));
end Behavioral;
