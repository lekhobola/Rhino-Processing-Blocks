--********************************************************************************
--* Company:        University of Cape Town									   
--* Engineer:       Lekhobola Joachim Tsoeunyane, lekhobola@gmail.com		       
--********************************************************************************
--* Create Date:    05-Jul-2014 22:07:35  				 										   
--* Design Name:    Pipelined R2^2 DIF-SDF FFT								       
--* Module Name:    fft1024_tf_rom_s0.vhd										   
--* Project Name:   RHINO SDR Processing Blocks								   
--* Target Devices: Xilinx - SPARTAN-6											   
--********************************************************************************
--* Dependencies: none															   
--********************************************************************************
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--********************************************************************************
--* This module implements the stage-0 of twiddle factor ROM for a 1024-point      
--* pipelined R2^2 DIF-SDF FFT. Each value is a complex number{imaginary,complex} 
--* ******************************************************************************
--* params:																	   
--*        addr_w - rom address bit width									       
--*        data_w - output data bit width										   
--* ports:																		   
--* 			[in]  addr	- Twidde factor ROM address to read					   
--* 			[out] doutr - Twiddle factor read from rom addr - real value	   
--* 			[out] douti - Twidder factor read from rom addr - imaginary value  
--********************************************************************************
--* Notes: Do not modify this file as it is auto-generated using matlab script    
--********************************************************************************
entity fft1024_tf_rom_s0 is
	generic(
		addr_w : natural := 10;
		data_w : natural := 16
	);
    port (
        addr  : in  std_logic_vector (addr_w - 1 downto 0);
        doutr : out std_logic_vector (data_w - 1 downto 0);
        douti : out  std_logic_vector(data_w - 1 downto 0)
 	);
end fft1024_tf_rom_s0;

architecture Behavioral of fft1024_tf_rom_s0 is
	type complex is array(0 to 1) of std_logic_vector(data_w - 1 downto 0);
	type rom_type is array(0 to (2 ** addr_w) - 1) of complex;

	constant rom : rom_type := (
								 ("0100000000000000","0000000000000000"),
								 ("0011111111111111","1111111100110111"),
								 ("0011111111111011","1111111001101110"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111101100","1111110011011100"),
								 ("0011111111100001","1111110000010011"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111111000100","1111101010000010"),
								 ("0011111110110001","1111100110111010"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111110000101","1111100000101010"),
								 ("0011111101101011","1111011101100011"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111100110000","1111010111010101"),
								 ("0011111100001111","1111010100001111"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111011000101","1111001110000100"),
								 ("0011111010011101","1111001010111111"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111001000101","1111000100110110"),
								 ("0011111000010101","1111000001110011"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110110101111","1110111011101110"),
								 ("0011110101111000","1110111000101101"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110100000011","1110110010101100"),
								 ("0011110011000101","1110101111101101"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110001000010","1110101001110000"),
								 ("0011101111111101","1110100110110100"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101101101101","1110100000111100"),
								 ("0011101100100001","1110011110000010"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101010000010","1110011000010001"),
								 ("0011101000110000","1110010101011001"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100110000100","1110001111101110"),
								 ("0011100100101011","1110001100111010"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100001110001","1110000111010101"),
								 ("0011100000010010","1110000100100100"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011101001011","1101111111000110"),
								 ("0011011011100101","1101111100011001"),
								 ("0011011001111101","1101111001101101"),
								 ("0011011000010010","1101110111000011"),
								 ("0011010110100101","1101110100011001"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010011000110","1101101111001011"),
								 ("0011010001010011","1101101100100110"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001101101000","1101100111100000"),
								 ("0011001011101111","1101100100111111"),
								 ("0011001001110100","1101100010100000"),
								 ("0011000111111000","1101100000000010"),
								 ("0011000101111001","1101011101100110"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000001110110","1101011000110010"),
								 ("0010111111110010","1101010110011011"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111011100100","1101010001110001"),
								 ("0010111001011010","1101001111011111"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110101000001","1101001010111111"),
								 ("0010110010110010","1101001000110001"),
								 ("0010110000100001","1101000110100110"),
								 ("0010101110001111","1101000100011100"),
								 ("0010101011111011","1101000010010100"),
								 ("0010101001100101","1101000000001110"),
								 ("0010100111001110","1100111110001010"),
								 ("0010100100110101","1100111100000111"),
								 ("0010100010011010","1100111010000111"),
								 ("0010011111111110","1100111000001000"),
								 ("0010011101100000","1100110110001100"),
								 ("0010011011000001","1100110100010001"),
								 ("0010011000100000","1100110010011000"),
								 ("0010010101111110","1100110000100001"),
								 ("0010010011011010","1100101110101101"),
								 ("0010010000110101","1100101100111010"),
								 ("0010001110001110","1100101011001001"),
								 ("0010001011100111","1100101001011011"),
								 ("0010001000111101","1100100111101110"),
								 ("0010000110010011","1100100110000011"),
								 ("0010000011100111","1100100100011011"),
								 ("0010000000111010","1100100010110101"),
								 ("0001111110001100","1100100001010000"),
								 ("0001111011011100","1100011111101110"),
								 ("0001111000101011","1100011110001111"),
								 ("0001110101111001","1100011100110001"),
								 ("0001110011000110","1100011011010101"),
								 ("0001110000010010","1100011001111100"),
								 ("0001101101011101","1100011000100101"),
								 ("0001101010100111","1100010111010000"),
								 ("0001100111101111","1100010101111110"),
								 ("0001100100110111","1100010100101101"),
								 ("0001100001111110","1100010011011111"),
								 ("0001011111000100","1100010010010011"),
								 ("0001011100001001","1100010001001010"),
								 ("0001011001001100","1100010000000011"),
								 ("0001010110010000","1100001110111110"),
								 ("0001010011010010","1100001101111011"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001101010100","1100001011111101"),
								 ("0001001010010100","1100001011000001"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000100010010","1100001001010001"),
								 ("0001000001010000","1100001000011101"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111011001010","1100000110111011"),
								 ("0000111000000110","1100000110001110"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110001111100","1100000100111011"),
								 ("0000101110110111","1100000100010101"),
								 ("0000101011110001","1100000011110001"),
								 ("0000101000101011","1100000011010000"),
								 ("0000100101100100","1100000010110001"),
								 ("0000100010011101","1100000010010101"),
								 ("0000011111010110","1100000001111011"),
								 ("0000011100001110","1100000001100100"),
								 ("0000011001000110","1100000001001111"),
								 ("0000010101111110","1100000000111100"),
								 ("0000010010110101","1100000000101100"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001100100100","1100000000010100"),
								 ("0000001001011011","1100000000001011"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000011001001","1100000000000001"),
								 ("0000000000000000","1100000000000000"),
								 ("1111111100110111","1100000000000001"),
								 ("1111111001101110","1100000000000101"),
								 ("1111110110100101","1100000000001011"),
								 ("1111110011011100","1100000000010100"),
								 ("1111110000010011","1100000000011111"),
								 ("1111101101001011","1100000000101100"),
								 ("1111101010000010","1100000000111100"),
								 ("1111100110111010","1100000001001111"),
								 ("1111100011110010","1100000001100100"),
								 ("1111100000101010","1100000001111011"),
								 ("1111011101100011","1100000010010101"),
								 ("1111011010011100","1100000010110001"),
								 ("1111010111010101","1100000011010000"),
								 ("1111010100001111","1100000011110001"),
								 ("1111010001001001","1100000100010101"),
								 ("1111001110000100","1100000100111011"),
								 ("1111001010111111","1100000101100011"),
								 ("1111000111111010","1100000110001110"),
								 ("1111000100110110","1100000110111011"),
								 ("1111000001110011","1100000111101011"),
								 ("1110111110110000","1100001000011101"),
								 ("1110111011101110","1100001001010001"),
								 ("1110111000101101","1100001010001000"),
								 ("1110110101101100","1100001011000001"),
								 ("1110110010101100","1100001011111101"),
								 ("1110101111101101","1100001100111011"),
								 ("1110101100101110","1100001101111011"),
								 ("1110101001110000","1100001110111110"),
								 ("1110100110110100","1100010000000011"),
								 ("1110100011110111","1100010001001010"),
								 ("1110100000111100","1100010010010011"),
								 ("1110011110000010","1100010011011111"),
								 ("1110011011001001","1100010100101101"),
								 ("1110011000010001","1100010101111110"),
								 ("1110010101011001","1100010111010000"),
								 ("1110010010100011","1100011000100101"),
								 ("1110001111101110","1100011001111100"),
								 ("1110001100111010","1100011011010101"),
								 ("1110001010000111","1100011100110001"),
								 ("1110000111010101","1100011110001111"),
								 ("1110000100100100","1100011111101110"),
								 ("1110000001110100","1100100001010000"),
								 ("1101111111000110","1100100010110101"),
								 ("1101111100011001","1100100100011011"),
								 ("1101111001101101","1100100110000011"),
								 ("1101110111000011","1100100111101110"),
								 ("1101110100011001","1100101001011011"),
								 ("1101110001110010","1100101011001001"),
								 ("1101101111001011","1100101100111010"),
								 ("1101101100100110","1100101110101101"),
								 ("1101101010000010","1100110000100001"),
								 ("1101100111100000","1100110010011000"),
								 ("1101100100111111","1100110100010001"),
								 ("1101100010100000","1100110110001100"),
								 ("1101100000000010","1100111000001000"),
								 ("1101011101100110","1100111010000111"),
								 ("1101011011001011","1100111100000111"),
								 ("1101011000110010","1100111110001010"),
								 ("1101010110011011","1101000000001110"),
								 ("1101010100000101","1101000010010100"),
								 ("1101010001110001","1101000100011100"),
								 ("1101001111011111","1101000110100110"),
								 ("1101001101001110","1101001000110001"),
								 ("1101001010111111","1101001010111111"),
								 ("1101001000110001","1101001101001110"),
								 ("1101000110100110","1101001111011111"),
								 ("1101000100011100","1101010001110001"),
								 ("1101000010010100","1101010100000101"),
								 ("1101000000001110","1101010110011011"),
								 ("1100111110001010","1101011000110010"),
								 ("1100111100000111","1101011011001011"),
								 ("1100111010000111","1101011101100110"),
								 ("1100111000001000","1101100000000010"),
								 ("1100110110001100","1101100010100000"),
								 ("1100110100010001","1101100100111111"),
								 ("1100110010011000","1101100111100000"),
								 ("1100110000100001","1101101010000010"),
								 ("1100101110101101","1101101100100110"),
								 ("1100101100111010","1101101111001011"),
								 ("1100101011001001","1101110001110010"),
								 ("1100101001011011","1101110100011001"),
								 ("1100100111101110","1101110111000011"),
								 ("1100100110000011","1101111001101101"),
								 ("1100100100011011","1101111100011001"),
								 ("1100100010110101","1101111111000110"),
								 ("1100100001010000","1110000001110100"),
								 ("1100011111101110","1110000100100100"),
								 ("1100011110001111","1110000111010101"),
								 ("1100011100110001","1110001010000111"),
								 ("1100011011010101","1110001100111010"),
								 ("1100011001111100","1110001111101110"),
								 ("1100011000100101","1110010010100011"),
								 ("1100010111010000","1110010101011001"),
								 ("1100010101111110","1110011000010001"),
								 ("1100010100101101","1110011011001001"),
								 ("1100010011011111","1110011110000010"),
								 ("1100010010010011","1110100000111100"),
								 ("1100010001001010","1110100011110111"),
								 ("1100010000000011","1110100110110100"),
								 ("1100001110111110","1110101001110000"),
								 ("1100001101111011","1110101100101110"),
								 ("1100001100111011","1110101111101101"),
								 ("1100001011111101","1110110010101100"),
								 ("1100001011000001","1110110101101100"),
								 ("1100001010001000","1110111000101101"),
								 ("1100001001010001","1110111011101110"),
								 ("1100001000011101","1110111110110000"),
								 ("1100000111101011","1111000001110011"),
								 ("1100000110111011","1111000100110110"),
								 ("1100000110001110","1111000111111010"),
								 ("1100000101100011","1111001010111111"),
								 ("1100000100111011","1111001110000100"),
								 ("1100000100010101","1111010001001001"),
								 ("1100000011110001","1111010100001111"),
								 ("1100000011010000","1111010111010101"),
								 ("1100000010110001","1111011010011100"),
								 ("1100000010010101","1111011101100011"),
								 ("1100000001111011","1111100000101010"),
								 ("1100000001100100","1111100011110010"),
								 ("1100000001001111","1111100110111010"),
								 ("1100000000111100","1111101010000010"),
								 ("1100000000101100","1111101101001011"),
								 ("1100000000011111","1111110000010011"),
								 ("1100000000010100","1111110011011100"),
								 ("1100000000001011","1111110110100101"),
								 ("1100000000000101","1111111001101110"),
								 ("1100000000000001","1111111100110111"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","1111111110011011"),
								 ("0011111111111111","1111111100110111"),
								 ("0011111111111101","1111111011010010"),
								 ("0011111111111011","1111111001101110"),
								 ("0011111111111000","1111111000001001"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111110001","1111110101000000"),
								 ("0011111111101100","1111110011011100"),
								 ("0011111111100111","1111110001111000"),
								 ("0011111111100001","1111110000010011"),
								 ("0011111111011011","1111101110101111"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111111001100","1111101011100110"),
								 ("0011111111000100","1111101010000010"),
								 ("0011111110111011","1111101000011110"),
								 ("0011111110110001","1111100110111010"),
								 ("0011111110100111","1111100101010110"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111110010001","1111100010001110"),
								 ("0011111110000101","1111100000101010"),
								 ("0011111101111000","1111011111000111"),
								 ("0011111101101011","1111011101100011"),
								 ("0011111101011101","1111011011111111"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111101000000","1111011000111001"),
								 ("0011111100110000","1111010111010101"),
								 ("0011111100100000","1111010101110010"),
								 ("0011111100001111","1111010100001111"),
								 ("0011111011111101","1111010010101100"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111011011000","1111001111100110"),
								 ("0011111011000101","1111001110000100"),
								 ("0011111010110001","1111001100100001"),
								 ("0011111010011101","1111001010111111"),
								 ("0011111010001000","1111001001011100"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111001011100","1111000110011000"),
								 ("0011111001000101","1111000100110110"),
								 ("0011111000101101","1111000011010101"),
								 ("0011111000010101","1111000001110011"),
								 ("0011110111111100","1111000000010010"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110111001001","1110111101001111"),
								 ("0011110110101111","1110111011101110"),
								 ("0011110110010011","1110111010001101"),
								 ("0011110101111000","1110111000101101"),
								 ("0011110101011011","1110110111001100"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110100100001","1110110100001100"),
								 ("0011110100000011","1110110010101100"),
								 ("0011110011100100","1110110001001100"),
								 ("0011110011000101","1110101111101101"),
								 ("0011110010100101","1110101110001101"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110001100100","1110101011001111"),
								 ("0011110001000010","1110101001110000"),
								 ("0011110000100000","1110101000010010"),
								 ("0011101111111101","1110100110110100"),
								 ("0011101111011010","1110100101010101"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101110010010","1110100010011010"),
								 ("0011101101101101","1110100000111100"),
								 ("0011101101000111","1110011111011111"),
								 ("0011101100100001","1110011110000010"),
								 ("0011101011111010","1110011100100101"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101010101011","1110011001101101"),
								 ("0011101010000010","1110011000010001"),
								 ("0011101001011001","1110010110110101"),
								 ("0011101000110000","1110010101011001"),
								 ("0011101000000110","1110010011111110"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100110110000","1110010001001000"),
								 ("0011100110000100","1110001111101110"),
								 ("0011100101011000","1110001110010100"),
								 ("0011100100101011","1110001100111010"),
								 ("0011100011111101","1110001011100000"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100010100001","1110001000101101"),
								 ("0011100001110001","1110000111010101"),
								 ("0011100001000010","1110000101111100"),
								 ("0011100000010010","1110000100100100"),
								 ("0011011111100001","1110000011001100"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011101111110","1110000000011101"),
								 ("0011011101001011","1101111111000110"),
								 ("0011011100011000","1101111101101111"),
								 ("0011011011100101","1101111100011001"),
								 ("0011011010110001","1101111011000011"),
								 ("0011011001111101","1101111001101101"),
								 ("0011011001001000","1101111000011000"),
								 ("0011011000010010","1101110111000011"),
								 ("0011010111011100","1101110101101110"),
								 ("0011010110100101","1101110100011001"),
								 ("0011010101101110","1101110011000101"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010011111111","1101110000011110"),
								 ("0011010011000110","1101101111001011"),
								 ("0011010010001101","1101101101111000"),
								 ("0011010001010011","1101101100100110"),
								 ("0011010000011001","1101101011010100"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001110100011","1101101000110001"),
								 ("0011001101101000","1101100111100000"),
								 ("0011001100101100","1101100110001111"),
								 ("0011001011101111","1101100100111111"),
								 ("0011001010110010","1101100011101111"),
								 ("0011001001110100","1101100010100000"),
								 ("0011001000110110","1101100001010001"),
								 ("0011000111111000","1101100000000010"),
								 ("0011000110111001","1101011110110100"),
								 ("0011000101111001","1101011101100110"),
								 ("0011000100111001","1101011100011001"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000010111000","1101011001111111"),
								 ("0011000001110110","1101011000110010"),
								 ("0011000000110100","1101010111100110"),
								 ("0010111111110010","1101010110011011"),
								 ("0010111110101111","1101010101010000"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111100101000","1101010010111011"),
								 ("0010111011100100","1101010001110001"),
								 ("0010111010011111","1101010000101000"),
								 ("0010111001011010","1101001111011111"),
								 ("0010111000010101","1101001110010110"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110110001000","1101001100000110"),
								 ("0010110101000001","1101001010111111"),
								 ("0010110011111010","1101001001111000"),
								 ("0010110010110010","1101001000110001"),
								 ("0010110001101010","1101000111101011"),
								 ("0010110000100001","1101000110100110"),
								 ("0010101111011000","1101000101100001"),
								 ("0010101110001111","1101000100011100"),
								 ("0010101101000101","1101000011011000"),
								 ("0010101011111011","1101000010010100"),
								 ("0010101010110000","1101000001010001"),
								 ("0010101001100101","1101000000001110"),
								 ("0010101000011010","1100111111001100"),
								 ("0010100111001110","1100111110001010"),
								 ("0010100110000001","1100111101001000"),
								 ("0010100100110101","1100111100000111"),
								 ("0010100011100111","1100111011000111"),
								 ("0010100010011010","1100111010000111"),
								 ("0010100001001100","1100111001000111"),
								 ("0010011111111110","1100111000001000"),
								 ("0010011110101111","1100110111001010"),
								 ("0010011101100000","1100110110001100"),
								 ("0010011100010001","1100110101001110"),
								 ("0010011011000001","1100110100010001"),
								 ("0010011001110001","1100110011010100"),
								 ("0010011000100000","1100110010011000"),
								 ("0010010111001111","1100110001011101"),
								 ("0010010101111110","1100110000100001"),
								 ("0010010100101100","1100101111100111"),
								 ("0010010011011010","1100101110101101"),
								 ("0010010010001000","1100101101110011"),
								 ("0010010000110101","1100101100111010"),
								 ("0010001111100010","1100101100000001"),
								 ("0010001110001110","1100101011001001"),
								 ("0010001100111011","1100101010010010"),
								 ("0010001011100111","1100101001011011"),
								 ("0010001010010010","1100101000100100"),
								 ("0010001000111101","1100100111101110"),
								 ("0010000111101000","1100100110111000"),
								 ("0010000110010011","1100100110000011"),
								 ("0010000100111101","1100100101001111"),
								 ("0010000011100111","1100100100011011"),
								 ("0010000010010001","1100100011101000"),
								 ("0010000000111010","1100100010110101"),
								 ("0001111111100011","1100100010000010"),
								 ("0001111110001100","1100100001010000"),
								 ("0001111100110100","1100100000011111"),
								 ("0001111011011100","1100011111101110"),
								 ("0001111010000100","1100011110111110"),
								 ("0001111000101011","1100011110001111"),
								 ("0001110111010011","1100011101011111"),
								 ("0001110101111001","1100011100110001"),
								 ("0001110100100000","1100011100000011"),
								 ("0001110011000110","1100011011010101"),
								 ("0001110001101100","1100011010101000"),
								 ("0001110000010010","1100011001111100"),
								 ("0001101110111000","1100011001010000"),
								 ("0001101101011101","1100011000100101"),
								 ("0001101100000010","1100010111111010"),
								 ("0001101010100111","1100010111010000"),
								 ("0001101001001011","1100010110100111"),
								 ("0001100111101111","1100010101111110"),
								 ("0001100110010011","1100010101010101"),
								 ("0001100100110111","1100010100101101"),
								 ("0001100011011011","1100010100000110"),
								 ("0001100001111110","1100010011011111"),
								 ("0001100000100001","1100010010111001"),
								 ("0001011111000100","1100010010010011"),
								 ("0001011101100110","1100010001101110"),
								 ("0001011100001001","1100010001001010"),
								 ("0001011010101011","1100010000100110"),
								 ("0001011001001100","1100010000000011"),
								 ("0001010111101110","1100001111100000"),
								 ("0001010110010000","1100001110111110"),
								 ("0001010100110001","1100001110011100"),
								 ("0001010011010010","1100001101111011"),
								 ("0001010001110011","1100001101011011"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001110110100","1100001100011100"),
								 ("0001001101010100","1100001011111101"),
								 ("0001001011110100","1100001011011111"),
								 ("0001001010010100","1100001011000001"),
								 ("0001001000110100","1100001010100101"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000101110011","1100001001101101"),
								 ("0001000100010010","1100001001010001"),
								 ("0001000010110001","1100001000110111"),
								 ("0001000001010000","1100001000011101"),
								 ("0000111111101110","1100001000000100"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111100101011","1100000111010011"),
								 ("0000111011001010","1100000110111011"),
								 ("0000111001101000","1100000110100100"),
								 ("0000111000000110","1100000110001110"),
								 ("0000110110100100","1100000101111000"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110011011111","1100000101001111"),
								 ("0000110001111100","1100000100111011"),
								 ("0000110000011010","1100000100101000"),
								 ("0000101110110111","1100000100010101"),
								 ("0000101101010100","1100000100000011"),
								 ("0000101011110001","1100000011110001"),
								 ("0000101010001110","1100000011100000"),
								 ("0000101000101011","1100000011010000"),
								 ("0000100111000111","1100000011000000"),
								 ("0000100101100100","1100000010110001"),
								 ("0000100100000001","1100000010100011"),
								 ("0000100010011101","1100000010010101"),
								 ("0000100000111001","1100000010001000"),
								 ("0000011111010110","1100000001111011"),
								 ("0000011101110010","1100000001101111"),
								 ("0000011100001110","1100000001100100"),
								 ("0000011010101010","1100000001011001"),
								 ("0000011001000110","1100000001001111"),
								 ("0000010111100010","1100000001000101"),
								 ("0000010101111110","1100000000111100"),
								 ("0000010100011010","1100000000110100"),
								 ("0000010010110101","1100000000101100"),
								 ("0000010001010001","1100000000100101"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001110001000","1100000000011001"),
								 ("0000001100100100","1100000000010100"),
								 ("0000001011000000","1100000000001111"),
								 ("0000001001011011","1100000000001011"),
								 ("0000000111110111","1100000000001000"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000100101110","1100000000000011"),
								 ("0000000011001001","1100000000000001"),
								 ("0000000001100101","1100000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0011111111111101","1111111011010010"),
								 ("0011111111110101","1111110110100101"),
								 ("0011111111100111","1111110001111000"),
								 ("0011111111010100","1111101101001011"),
								 ("0011111110111011","1111101000011110"),
								 ("0011111110011100","1111100011110010"),
								 ("0011111101111000","1111011111000111"),
								 ("0011111101001111","1111011010011100"),
								 ("0011111100100000","1111010101110010"),
								 ("0011111011101011","1111010001001001"),
								 ("0011111010110001","1111001100100001"),
								 ("0011111001110010","1111000111111010"),
								 ("0011111000101101","1111000011010101"),
								 ("0011110111100011","1110111110110000"),
								 ("0011110110010011","1110111010001101"),
								 ("0011110100111111","1110110101101100"),
								 ("0011110011100100","1110110001001100"),
								 ("0011110010000101","1110101100101110"),
								 ("0011110000100000","1110101000010010"),
								 ("0011101110110110","1110100011110111"),
								 ("0011101101000111","1110011111011111"),
								 ("0011101011010011","1110011011001001"),
								 ("0011101001011001","1110010110110101"),
								 ("0011100111011011","1110010010100011"),
								 ("0011100101011000","1110001110010100"),
								 ("0011100011001111","1110001010000111"),
								 ("0011100001000010","1110000101111100"),
								 ("0011011110110000","1110000001110100"),
								 ("0011011100011000","1101111101101111"),
								 ("0011011001111101","1101111001101101"),
								 ("0011010111011100","1101110101101110"),
								 ("0011010100110111","1101110001110010"),
								 ("0011010010001101","1101101101111000"),
								 ("0011001111011111","1101101010000010"),
								 ("0011001100101100","1101100110001111"),
								 ("0011001001110100","1101100010100000"),
								 ("0011000110111001","1101011110110100"),
								 ("0011000011111001","1101011011001011"),
								 ("0011000000110100","1101010111100110"),
								 ("0010111101101100","1101010100000101"),
								 ("0010111010011111","1101010000101000"),
								 ("0010110111001111","1101001101001110"),
								 ("0010110011111010","1101001001111000"),
								 ("0010110000100001","1101000110100110"),
								 ("0010101101000101","1101000011011000"),
								 ("0010101001100101","1101000000001110"),
								 ("0010100110000001","1100111101001000"),
								 ("0010100010011010","1100111010000111"),
								 ("0010011110101111","1100110111001010"),
								 ("0010011011000001","1100110100010001"),
								 ("0010010111001111","1100110001011101"),
								 ("0010010011011010","1100101110101101"),
								 ("0010001111100010","1100101100000001"),
								 ("0010001011100111","1100101001011011"),
								 ("0010000111101000","1100100110111000"),
								 ("0010000011100111","1100100100011011"),
								 ("0001111111100011","1100100010000010"),
								 ("0001111011011100","1100011111101110"),
								 ("0001110111010011","1100011101011111"),
								 ("0001110011000110","1100011011010101"),
								 ("0001101110111000","1100011001010000"),
								 ("0001101010100111","1100010111010000"),
								 ("0001100110010011","1100010101010101"),
								 ("0001100001111110","1100010011011111"),
								 ("0001011101100110","1100010001101110"),
								 ("0001011001001100","1100010000000011"),
								 ("0001010100110001","1100001110011100"),
								 ("0001010000010011","1100001100111011"),
								 ("0001001011110100","1100001011011111"),
								 ("0001000111010011","1100001010001000"),
								 ("0001000010110001","1100001000110111"),
								 ("0000111110001101","1100000111101011"),
								 ("0000111001101000","1100000110100100"),
								 ("0000110101000001","1100000101100011"),
								 ("0000110000011010","1100000100101000"),
								 ("0000101011110001","1100000011110001"),
								 ("0000100111000111","1100000011000000"),
								 ("0000100010011101","1100000010010101"),
								 ("0000011101110010","1100000001101111"),
								 ("0000011001000110","1100000001001111"),
								 ("0000010100011010","1100000000110100"),
								 ("0000001111101101","1100000000011111"),
								 ("0000001011000000","1100000000001111"),
								 ("0000000110010010","1100000000000101"),
								 ("0000000001100101","1100000000000000"),
								 ("1111111100110111","1100000000000001"),
								 ("1111111000001001","1100000000001000"),
								 ("1111110011011100","1100000000010100"),
								 ("1111101110101111","1100000000100101"),
								 ("1111101010000010","1100000000111100"),
								 ("1111100101010110","1100000001011001"),
								 ("1111100000101010","1100000001111011"),
								 ("1111011011111111","1100000010100011"),
								 ("1111010111010101","1100000011010000"),
								 ("1111010010101100","1100000100000011"),
								 ("1111001110000100","1100000100111011"),
								 ("1111001001011100","1100000101111000"),
								 ("1111000100110110","1100000110111011"),
								 ("1111000000010010","1100001000000100"),
								 ("1110111011101110","1100001001010001"),
								 ("1110110111001100","1100001010100101"),
								 ("1110110010101100","1100001011111101"),
								 ("1110101110001101","1100001101011011"),
								 ("1110101001110000","1100001110111110"),
								 ("1110100101010101","1100010000100110"),
								 ("1110100000111100","1100010010010011"),
								 ("1110011100100101","1100010100000110"),
								 ("1110011000010001","1100010101111110"),
								 ("1110010011111110","1100010111111010"),
								 ("1110001111101110","1100011001111100"),
								 ("1110001011100000","1100011100000011"),
								 ("1110000111010101","1100011110001111"),
								 ("1110000011001100","1100100000011111"),
								 ("1101111111000110","1100100010110101"),
								 ("1101111011000011","1100100101001111"),
								 ("1101110111000011","1100100111101110"),
								 ("1101110011000101","1100101010010010"),
								 ("1101101111001011","1100101100111010"),
								 ("1101101011010100","1100101111100111"),
								 ("1101100111100000","1100110010011000"),
								 ("1101100011101111","1100110101001110"),
								 ("1101100000000010","1100111000001000"),
								 ("1101011100011001","1100111011000111"),
								 ("1101011000110010","1100111110001010"),
								 ("1101010101010000","1101000001010001"),
								 ("1101010001110001","1101000100011100"),
								 ("1101001110010110","1101000111101011"),
								 ("1101001010111111","1101001010111111"),
								 ("1101000111101011","1101001110010110"),
								 ("1101000100011100","1101010001110001"),
								 ("1101000001010001","1101010101010000"),
								 ("1100111110001010","1101011000110010"),
								 ("1100111011000111","1101011100011001"),
								 ("1100111000001000","1101100000000010"),
								 ("1100110101001110","1101100011101111"),
								 ("1100110010011000","1101100111100000"),
								 ("1100101111100111","1101101011010100"),
								 ("1100101100111010","1101101111001011"),
								 ("1100101010010010","1101110011000101"),
								 ("1100100111101110","1101110111000011"),
								 ("1100100101001111","1101111011000011"),
								 ("1100100010110101","1101111111000110"),
								 ("1100100000011111","1110000011001100"),
								 ("1100011110001111","1110000111010101"),
								 ("1100011100000011","1110001011100000"),
								 ("1100011001111100","1110001111101110"),
								 ("1100010111111010","1110010011111110"),
								 ("1100010101111110","1110011000010001"),
								 ("1100010100000110","1110011100100101"),
								 ("1100010010010011","1110100000111100"),
								 ("1100010000100110","1110100101010101"),
								 ("1100001110111110","1110101001110000"),
								 ("1100001101011011","1110101110001101"),
								 ("1100001011111101","1110110010101100"),
								 ("1100001010100101","1110110111001100"),
								 ("1100001001010001","1110111011101110"),
								 ("1100001000000100","1111000000010010"),
								 ("1100000110111011","1111000100110110"),
								 ("1100000101111000","1111001001011100"),
								 ("1100000100111011","1111001110000100"),
								 ("1100000100000011","1111010010101100"),
								 ("1100000011010000","1111010111010101"),
								 ("1100000010100011","1111011011111111"),
								 ("1100000001111011","1111100000101010"),
								 ("1100000001011001","1111100101010110"),
								 ("1100000000111100","1111101010000010"),
								 ("1100000000100101","1111101110101111"),
								 ("1100000000010100","1111110011011100"),
								 ("1100000000001000","1111111000001001"),
								 ("1100000000000001","1111111100110111"),
								 ("1100000000000000","0000000001100101"),
								 ("1100000000000101","0000000110010010"),
								 ("1100000000001111","0000001011000000"),
								 ("1100000000011111","0000001111101101"),
								 ("1100000000110100","0000010100011010"),
								 ("1100000001001111","0000011001000110"),
								 ("1100000001101111","0000011101110010"),
								 ("1100000010010101","0000100010011101"),
								 ("1100000011000000","0000100111000111"),
								 ("1100000011110001","0000101011110001"),
								 ("1100000100101000","0000110000011010"),
								 ("1100000101100011","0000110101000001"),
								 ("1100000110100100","0000111001101000"),
								 ("1100000111101011","0000111110001101"),
								 ("1100001000110111","0001000010110001"),
								 ("1100001010001000","0001000111010011"),
								 ("1100001011011111","0001001011110100"),
								 ("1100001100111011","0001010000010011"),
								 ("1100001110011100","0001010100110001"),
								 ("1100010000000011","0001011001001100"),
								 ("1100010001101110","0001011101100110"),
								 ("1100010011011111","0001100001111110"),
								 ("1100010101010101","0001100110010011"),
								 ("1100010111010000","0001101010100111"),
								 ("1100011001010000","0001101110111000"),
								 ("1100011011010101","0001110011000110"),
								 ("1100011101011111","0001110111010011"),
								 ("1100011111101110","0001111011011100"),
								 ("1100100010000010","0001111111100011"),
								 ("1100100100011011","0010000011100111"),
								 ("1100100110111000","0010000111101000"),
								 ("1100101001011011","0010001011100111"),
								 ("1100101100000001","0010001111100010"),
								 ("1100101110101101","0010010011011010"),
								 ("1100110001011101","0010010111001111"),
								 ("1100110100010001","0010011011000001"),
								 ("1100110111001010","0010011110101111"),
								 ("1100111010000111","0010100010011010"),
								 ("1100111101001000","0010100110000001"),
								 ("1101000000001110","0010101001100101"),
								 ("1101000011011000","0010101101000101"),
								 ("1101000110100110","0010110000100001"),
								 ("1101001001111000","0010110011111010"),
								 ("1101001101001110","0010110111001111"),
								 ("1101010000101000","0010111010011111"),
								 ("1101010100000101","0010111101101100"),
								 ("1101010111100110","0011000000110100"),
								 ("1101011011001011","0011000011111001"),
								 ("1101011110110100","0011000110111001"),
								 ("1101100010100000","0011001001110100"),
								 ("1101100110001111","0011001100101100"),
								 ("1101101010000010","0011001111011111"),
								 ("1101101101111000","0011010010001101"),
								 ("1101110001110010","0011010100110111"),
								 ("1101110101101110","0011010111011100"),
								 ("1101111001101101","0011011001111101"),
								 ("1101111101101111","0011011100011000"),
								 ("1110000001110100","0011011110110000"),
								 ("1110000101111100","0011100001000010"),
								 ("1110001010000111","0011100011001111"),
								 ("1110001110010100","0011100101011000"),
								 ("1110010010100011","0011100111011011"),
								 ("1110010110110101","0011101001011001"),
								 ("1110011011001001","0011101011010011"),
								 ("1110011111011111","0011101101000111"),
								 ("1110100011110111","0011101110110110"),
								 ("1110101000010010","0011110000100000"),
								 ("1110101100101110","0011110010000101"),
								 ("1110110001001100","0011110011100100"),
								 ("1110110101101100","0011110100111111"),
								 ("1110111010001101","0011110110010011"),
								 ("1110111110110000","0011110111100011"),
								 ("1111000011010101","0011111000101101"),
								 ("1111000111111010","0011111001110010"),
								 ("1111001100100001","0011111010110001"),
								 ("1111010001001001","0011111011101011"),
								 ("1111010101110010","0011111100100000"),
								 ("1111011010011100","0011111101001111"),
								 ("1111011111000111","0011111101111000"),
								 ("1111100011110010","0011111110011100"),
								 ("1111101000011110","0011111110111011"),
								 ("1111101101001011","0011111111010100"),
								 ("1111110001111000","0011111111100111"),
								 ("1111110110100101","0011111111110101"),
								 ("1111111011010010","0011111111111101"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000"),
								 ("0100000000000000","0000000000000000")
							   );
begin
	doutr <= std_logic_vector(rom(conv_integer(addr))(0));
	douti <= std_logic_vector(rom(conv_integer(addr))(1));
end Behavioral;
